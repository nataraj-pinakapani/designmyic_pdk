magic
tech sky130A
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__dfl1sd__example_55959141808123  sky130_fd_pr__dfl1sd__example_55959141808123_0
timestamp 1663361622
transform -1 0 -14 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808123  sky130_fd_pr__dfl1sd__example_55959141808123_1
timestamp 1663361622
transform 1 0 800 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 32319282
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 32318168
<< end >>
