/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos/begin_of_life/worst.spice