magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 32 163 52 167 6 G_PAD
port 3 nsew signal bidirectional
rlabel � s 21 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 21 0 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 21 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 21 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 21 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 21 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 21 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 21 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 2 54 2 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 2 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 20 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 3 54 3 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 3 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 19 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 4 54 4 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 4 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 5 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel � s 18 5 54 10 6 BDY2_B2B
port 4 nsew ground bidirectional
rlabel 
 s 54 164 60 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 100 60 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 100 60 100 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 100 60 100 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 165 60 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 100 60 100 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 165 60 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 100 60 100 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 165 60 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 99 60 100 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 165 60 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 99 60 99 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 165 60 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 54 99 60 99 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 165 60 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 99 60 99 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 166 60 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 99 60 99 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 166 60 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 99 60 99 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 166 60 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 99 60 99 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 166 60 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 98 60 99 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 166 60 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 98 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 53 166 60 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 98 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 166 60 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 98 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 167 60 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 98 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 167 60 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 98 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 167 60 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 98 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 98 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 167 60 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 97 60 98 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 167 60 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 52 97 60 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 167 60 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 97 60 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 167 60 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 97 60 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 168 60 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 97 59 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 168 60 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 97 59 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 168 60 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 96 59 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 168 60 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 96 59 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 51 168 60 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 96 59 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 168 60 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 96 59 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 169 60 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 96 59 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 169 60 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 96 58 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 169 60 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 96 58 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 169 60 190 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 95 58 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 50 95 58 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 49 95 58 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 49 95 58 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 49 95 57 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 49 95 57 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 49 95 57 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 49 94 57 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 49 94 57 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 48 94 57 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 48 94 57 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 48 94 56 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 48 94 56 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 48 93 56 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 48 93 56 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 47 93 56 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 47 93 56 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 47 93 56 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 47 93 55 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 47 93 55 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 47 92 55 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 47 92 55 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 46 92 55 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 46 92 55 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 46 92 54 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 46 92 54 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 46 92 54 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 46 91 54 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 46 91 54 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 45 91 54 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 45 91 54 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 45 91 53 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 45 91 53 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 45 90 53 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 45 90 53 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 44 90 53 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 44 90 53 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 44 90 53 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 44 90 52 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 44 90 52 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 44 89 52 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 44 89 52 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 89 52 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 89 52 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 89 51 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 89 51 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 89 51 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 164 49 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 97 49 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 97 49 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 97 49 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 96 48 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 96 48 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 96 48 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 96 48 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 96 48 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 96 48 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 96 48 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 95 47 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 95 47 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 95 47 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 88 51 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 164 49 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 95 47 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 88 51 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 164 49 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 43 88 51 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 95 47 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 165 49 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 88 51 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 95 47 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 165 49 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 88 51 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 95 47 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 165 49 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 88 51 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 94 46 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 165 49 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 88 51 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 94 46 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 165 49 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 87 51 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 94 46 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 165 49 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 87 51 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 87 51 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 87 51 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 87 51 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 86 51 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 86 50 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 86 50 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 86 50 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 86 50 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 86 50 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 86 50 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 85 49 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 85 49 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 85 49 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 85 49 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 85 49 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 85 49 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 85 49 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 94 46 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 42 84 49 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 165 49 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 94 46 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 84 49 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 166 49 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 94 46 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 84 49 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 166 49 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 94 46 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 84 49 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 166 49 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 93 45 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 166 49 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 93 45 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 166 49 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 93 45 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 41 166 49 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 93 45 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 167 49 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 93 45 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 167 49 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 93 45 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 167 49 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 92 45 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 167 49 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 92 44 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 167 49 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 92 44 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 167 49 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 92 44 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 40 167 49 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 92 44 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 168 49 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 92 44 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 168 49 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 92 44 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 168 49 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 91 43 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 168 49 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 91 43 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 168 49 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 91 43 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 168 49 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 39 91 43 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 168 49 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 91 43 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 169 49 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 91 43 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 169 49 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 91 43 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 169 49 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 169 49 190 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 90 42 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 35 86 39 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 35 85 39 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 35 85 39 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 84 39 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 86 39 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 84 40 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 86 39 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 84 40 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 86 39 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 84 40 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 87 39 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 87 39 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 34 87 39 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 33 87 39 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 33 87 39 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 33 87 39 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 33 88 40 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 33 88 40 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 33 88 40 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 33 88 40 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 32 88 40 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 32 88 40 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 32 88 40 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 32 89 41 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 32 89 41 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 32 89 41 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 32 89 41 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 31 89 41 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 31 89 41 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 31 89 41 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 31 90 42 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 31 90 42 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 31 90 42 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 90 42 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 90 42 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 90 42 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 90 35 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 91 35 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 91 35 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 91 34 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 30 91 34 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 29 91 34 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 29 91 34 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 29 91 34 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 29 92 34 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 29 92 34 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 29 92 33 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 29 92 33 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 28 92 33 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 28 92 33 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 28 92 33 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 28 93 33 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 28 93 33 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 28 93 32 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 93 32 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 93 32 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 93 32 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 93 32 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 94 32 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 94 32 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 94 32 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 27 94 32 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 94 32 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 94 32 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 94 32 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 167 37 190 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 167 37 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 167 37 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 167 37 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 167 36 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 167 36 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 167 36 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 166 36 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 166 36 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 166 36 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 166 35 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 166 35 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 166 35 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 166 35 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 165 35 166 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 165 35 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 165 35 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 165 34 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 165 34 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 165 34 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 165 34 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 164 34 165 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 164 34 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 164 34 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 164 33 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 164 33 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 164 33 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 163 33 164 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 163 33 163 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 163 33 163 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 163 32 163 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 163 32 163 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 163 32 163 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 163 32 163 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 95 32 163 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 83 49 83 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 77 49 83 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 77 49 77 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 77 49 77 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 76 48 77 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 76 48 76 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 76 48 76 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 76 48 76 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 76 48 76 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 76 48 76 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 48 76 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 47 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 47 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 47 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 47 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 47 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 40 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 75 40 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 74 40 75 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 74 40 74 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 74 40 74 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 74 40 74 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 74 40 74 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 74 39 74 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 74 39 74 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 73 39 74 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 73 39 73 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 73 39 73 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 73 39 73 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 73 39 73 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 73 38 73 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 72 38 73 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 72 38 72 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 72 38 72 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 72 38 72 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 72 38 72 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 72 37 72 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 72 37 72 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 71 37 72 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 71 37 71 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 71 37 71 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 0 37 71 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 83 49 83 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 83 49 83 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 26 83 49 83 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 25 83 49 83 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 25 83 49 83 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 25 83 49 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 25 84 49 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 25 84 49 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 25 84 49 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 25 84 33 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 84 33 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 84 32 84 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 84 32 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 85 32 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 86 32 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 85 32 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 85 32 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 85 32 85 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 86 32 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 86 32 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 86 32 86 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 24 86 32 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 23 87 32 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 23 87 32 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 23 87 31 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 23 87 31 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 23 87 31 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 23 87 31 87 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 22 87 31 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 22 88 31 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 22 88 30 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 22 88 30 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 22 88 30 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 22 88 30 88 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 22 88 30 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 21 89 30 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 21 89 30 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 21 89 29 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 21 89 29 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 21 89 29 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 21 89 29 89 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 21 89 29 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 20 90 29 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 20 90 29 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 20 90 28 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 20 90 28 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 20 90 28 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 20 90 28 90 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 19 90 28 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 19 91 28 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 19 91 27 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 19 91 27 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 19 91 27 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 19 91 27 91 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 19 91 27 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 18 92 27 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 18 92 27 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 18 92 26 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 18 92 26 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 18 92 26 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 18 92 26 92 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 18 92 26 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 17 93 26 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 17 93 26 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 17 93 25 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 17 93 25 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 17 93 25 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 17 93 25 93 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 93 25 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 94 25 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 94 24 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 94 24 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 94 24 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 94 24 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 171 25 190 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 171 25 171 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 170 25 171 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 170 25 170 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 170 25 170 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 170 24 170 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 170 24 170 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 170 24 170 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 170 24 170 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 169 24 170 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 169 24 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 169 24 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 169 23 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 169 23 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 169 23 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 168 23 169 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 168 23 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 168 23 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 168 23 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 168 22 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 168 22 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 168 22 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 167 22 168 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 167 22 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 167 22 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 97 22 167 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 97 22 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 97 22 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 96 22 97 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 96 22 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 96 22 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 96 22 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 96 22 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 96 23 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 96 23 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 95 23 96 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 95 23 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 95 23 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 95 23 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 95 23 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 95 24 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 94 24 95 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 16 94 24 94 6 DRN_LVC1
port 5 nsew power bidirectional
rlabel 
 s 38 0 49 69 6 DRN_LVC2
port 6 nsew power bidirectional
rlabel 
 s 1 94 13 171 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 94 13 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 94 13 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 94 13 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 94 13 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 94 13 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 93 14 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 93 14 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 93 14 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 93 14 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 93 14 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 93 14 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 93 14 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 92 15 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 92 15 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 92 15 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 92 15 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 92 15 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 92 15 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 92 16 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 91 16 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 91 16 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 91 16 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 91 16 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 91 16 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 91 16 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 90 17 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 90 17 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 90 17 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 90 17 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 90 17 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 90 17 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 90 17 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 89 18 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 89 18 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 89 18 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 89 18 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 89 18 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 89 18 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 89 19 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 88 19 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 88 19 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 88 19 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 88 19 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 88 19 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 88 19 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 87 20 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 87 20 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 87 20 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 87 20 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 87 20 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 87 20 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 87 20 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 86 21 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 86 21 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 86 21 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 86 21 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 86 21 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 86 21 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 86 22 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 85 22 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 85 22 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 85 22 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 85 22 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 85 22 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 85 22 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 84 23 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 84 23 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 84 23 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 84 23 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 84 23 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 84 23 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 84 23 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 83 24 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 83 24 83 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 83 24 83 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 83 24 83 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 83 24 83 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 83 24 83 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 1 0 25 83 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 62 96 75 172 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 62 96 75 96 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 62 96 75 96 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 62 95 75 96 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 62 95 75 95 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 62 95 75 95 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 61 95 75 95 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 61 95 75 95 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 61 95 75 95 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 61 95 75 95 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 61 94 75 95 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 61 94 75 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 61 94 75 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 60 94 75 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 60 94 75 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 60 94 75 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 60 93 75 94 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 60 93 75 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 60 93 75 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 59 93 75 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 59 93 75 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 59 93 75 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 59 93 75 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 59 92 75 93 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 59 92 75 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 59 92 75 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 58 92 75 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 58 92 75 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 58 92 75 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 58 92 75 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 58 91 75 92 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 58 91 75 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 58 91 75 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 57 91 75 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 57 91 75 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 57 91 75 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 57 90 75 91 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 57 90 75 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 57 90 75 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 56 90 75 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 56 90 75 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 56 90 75 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 56 90 75 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 56 89 75 90 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 56 89 75 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 56 89 75 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 55 89 75 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 55 89 75 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 55 89 75 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 55 89 75 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 55 88 75 89 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 55 88 75 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 55 88 75 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 54 88 75 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 54 88 75 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 54 88 75 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 54 87 75 88 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 54 87 75 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 54 87 75 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 53 87 75 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 53 87 75 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 53 87 75 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 53 87 75 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 53 86 75 87 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 53 86 75 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 53 86 75 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 52 86 75 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 52 86 75 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 52 86 75 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 52 86 75 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 52 85 75 86 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 52 85 75 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 52 85 75 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 51 85 75 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 51 85 75 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 51 85 75 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 51 84 75 85 6 G_CORE
port 7 nsew ground bidirectional
rlabel 
 s 51 0 75 84 6 G_CORE
port 7 nsew ground bidirectional
rlabel  s 26 0 28 0 8 OGC_LVC
port 8 nsew power bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 9 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 9 17 9 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 8 17 9 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 8 17 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 8 17 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 8 17 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 17 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 8 17 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 18 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 56 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 8 17 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 56 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 8 17 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 12 10 56 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 68 194 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 15 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 15 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 15 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 15 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 15 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 15 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 191 15 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 191 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 185 14 190 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 14 185 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 14 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 14 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 14 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 14 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 14 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 68 184 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 15 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 15 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 15 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 15 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 15 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 15 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 181 15 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 181 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 180 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 175 14 180 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 175 14 175 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 175 14 175 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 14 175 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 14 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 14 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 14 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 14 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 14 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 15 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 15 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 15 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 15 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 15 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 15 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 174 15 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 68 174 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 171 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 165 14 170 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 165 14 165 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 165 14 165 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 14 165 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 14 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 14 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 14 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 14 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 14 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 15 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 15 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 15 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 15 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 15 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 15 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 164 15 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 68 164 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 161 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 160 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 155 14 160 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 155 14 155 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 155 14 155 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 14 155 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 14 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 14 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 14 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 14 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 14 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 15 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 15 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 15 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 15 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 15 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 15 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 154 15 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 68 154 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 15 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 15 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 15 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 15 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 15 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 15 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 151 15 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 151 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 150 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 145 14 150 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 145 14 145 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 145 14 145 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 14 145 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 14 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 14 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 14 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 14 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 14 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 15 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 15 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 15 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 15 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 15 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 15 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 144 15 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 68 144 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 15 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 15 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 15 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 15 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 15 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 15 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 141 15 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 141 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 140 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 135 14 140 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 135 14 135 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 135 14 135 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 14 135 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 14 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 14 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 14 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 14 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 14 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 15 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 15 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 15 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 15 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 15 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 15 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 134 15 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 131 68 134 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 131 15 131 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 131 15 131 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 131 15 131 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 131 15 131 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 131 15 131 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 131 15 131 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 15 131 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 130 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 75 14 130 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 74 14 75 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 74 14 74 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 74 14 74 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 74 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 25 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 14 25 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 24 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 15 24 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 15 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 23 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 16 23 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 16 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 22 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 17 22 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 17 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 21 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 18 21 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 18 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 20 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 19 20 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 19 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 19 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 20 19 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 20 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 18 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 17 21 18 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 17 22 17 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 17 22 17 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 17 22 17 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 17 22 17 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 17 22 17 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 10 56 17 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 10 11 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 10 11 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 10 11 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 10 11 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 10 10 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 10 10 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 8 10 10 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 8 10 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 8 10 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 8 11 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 8 11 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 8 11 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 8 11 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 8 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 5 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 17 5 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 17 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 4 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 18 4 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 3 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 19 3 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 2 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 1 20 2 6 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 1 0 20 1 8 SRC_BDY_LVC1
port 9 nsew ground bidirectional
rlabel � s 66 74 68 99 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 45 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 45 75 45 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 35 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 35 75 35 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 65 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 65 75 65 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 55 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 55 75 55 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 55 75 55 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 45 75 45 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 35 75 35 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 65 75 65 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 54 75 55 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 44 75 45 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 34 75 35 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 64 75 65 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 50 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 70 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 60 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 74 68 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 50 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 40 75 40 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 30 75 30 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 70 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 66 60 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 74 69 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 40 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 30 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 71 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 61 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 74 69 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 41 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 71 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 61 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 74 69 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 41 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 71 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 61 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 74 69 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 41 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 71 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 61 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 25 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 41 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 71 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 61 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 25 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 41 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 71 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 61 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 54 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 44 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 34 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 41 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 71 75 71 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 64 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 61 75 61 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 51 75 51 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 41 75 41 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 31 75 31 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 65 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 24 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 24 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 64 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 23 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 23 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 63 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 62 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 62 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 62 22 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 10 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 10 75 10 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 10 75 10 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 10 75 10 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 10 75 10 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 10 75 10 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 10 75 10 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 9 75 10 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 18 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 18 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 56 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 9 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 8 75 9 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 19 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 19 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 20 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 55 20 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 20 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 20 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 20 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 20 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 8 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 20 75 20 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 20 75 22 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 54 0 75 8 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 16 71 75 74 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 16 61 75 64 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 16 51 75 54 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 16 41 75 44 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel � s 16 31 75 34 6 SRC_BDY_LVC2
port 10 nsew ground bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 11 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 11 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 11 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 11 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 12 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 12 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 12 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 12 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 13 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 13 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 13 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 13 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 15 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 15 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 15 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 15 nsew power bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 16 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 16 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 16 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 16 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 16 nsew ground bidirectional
rlabel  s 74 46 75 46 6 VSSA
port 16 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 16 nsew ground bidirectional
rlabel  s 74 54 75 55 6 VSSA
port 16 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 16 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 16 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 16 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 16 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 17 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 17 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 17 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 17 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 18 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 18 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 18 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 18 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 18 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 18 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 18 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 18 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 19 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 19 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 19 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 19 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 20 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 20 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 20 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 20 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 198
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
