magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< metal4 >>
rect 0 34750 1000 39593
rect 0 13600 1000 18593
rect 0 12410 1000 13300
rect 0 11240 1000 12130
rect 0 10218 1000 10814
rect 0 9266 1000 9862
rect 0 7910 1000 8840
rect 0 5970 1000 6660
rect 0 4760 1000 5690
rect 0 3550 1000 4480
rect 0 1370 1000 2300
rect 0 0 1000 1090
<< metal5 >>
rect 0 34750 1000 39593
rect 0 13600 1000 18590
rect 0 12430 1000 13280
rect 0 11260 1000 12110
rect 0 7930 1000 8820
rect 0 5990 1000 6640
rect 0 4780 1000 5670
rect 0 3570 1000 4460
rect 0 1390 1000 2280
rect 0 20 1000 1070
<< labels >>
flabel metal4 s 800 10218 1000 10814 0 FreeSans 1000 0 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 0 10218 200 10814 0 FreeSans 1000 0 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 800 9266 1000 9862 0 FreeSans 1000 0 0 0 AMUXBUS_B
port 2 nsew
flabel metal4 s 0 9266 200 9862 0 FreeSans 1000 0 0 0 AMUXBUS_B
port 2 nsew
flabel metal5 s 0 5990 200 6640 0 FreeSans 1000 0 0 0 VSWITCH
port 3 nsew
flabel metal4 s 0 5970 200 6660 0 FreeSans 1000 0 0 0 VSWITCH
port 3 nsew
flabel metal5 s 800 5990 1000 6640 0 FreeSans 1000 0 0 0 VSWITCH
port 3 nsew
flabel metal4 s 800 5970 1000 6660 0 FreeSans 1000 0 0 0 VSWITCH
port 3 nsew
flabel metal5 s 0 12430 200 13280 0 FreeSans 1000 0 0 0 VDDIO_Q
port 4 nsew
flabel metal5 s 800 12430 1000 13280 0 FreeSans 1000 0 0 0 VDDIO_Q
port 4 nsew
flabel metal4 s 800 12410 1000 13300 0 FreeSans 1000 0 0 0 VDDIO_Q
port 4 nsew
flabel metal5 s 0 20 200 1070 0 FreeSans 1000 0 0 0 VCCHIB
port 5 nsew
flabel metal4 s 0 0 200 1090 0 FreeSans 1000 0 0 0 VCCHIB
port 5 nsew
flabel metal5 s 800 20 1000 1070 0 FreeSans 1000 0 0 0 VCCHIB
port 5 nsew
flabel metal4 s 800 0 1000 1090 0 FreeSans 1000 0 0 0 VCCHIB
port 5 nsew
rlabel metal4 s 800 3550 1000 4480 4 VDDIO
port 6 nsew
flabel metal5 s 0 13600 200 18590 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal4 s 0 13600 200 18593 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal5 s 0 3570 200 4460 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal4 s 0 3550 200 4480 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal5 s 800 13600 1000 18590 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal4 s 800 13600 1000 18593 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal5 s 800 3570 1000 4460 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal4 s 900 4015 900 4015 0 FreeSans 1000 0 0 0 VDDIO
port 6 nsew
flabel metal5 s 0 1390 200 2280 0 FreeSans 1000 0 0 0 VCCD
port 7 nsew
flabel metal4 s 0 1370 200 2300 0 FreeSans 1000 0 0 0 VCCD
port 7 nsew
flabel metal5 s 800 1390 1000 2280 0 FreeSans 1000 0 0 0 VCCD
port 7 nsew
flabel metal4 s 800 1370 1000 2300 0 FreeSans 1000 0 0 0 VCCD
port 7 nsew
flabel metal5 s 0 4780 200 5670 0 FreeSans 1000 0 0 0 VSSIO
port 8 nsew
flabel metal4 s 0 4760 200 5690 0 FreeSans 1000 0 0 0 VSSIO
port 8 nsew
flabel metal5 s 0 34750 200 39593 0 FreeSans 1000 0 0 0 VSSIO
port 8 nsew
flabel metal5 s 800 4780 1000 5670 0 FreeSans 1000 0 0 0 VSSIO
port 8 nsew
flabel metal4 s 800 4760 1000 5690 0 FreeSans 1000 0 0 0 VSSIO
port 8 nsew
flabel metal5 s 800 34750 1000 39593 0 FreeSans 1000 0 0 0 VSSIO
port 8 nsew
flabel metal5 s 0 7930 200 8820 0 FreeSans 1000 0 0 0 VSSD
port 9 nsew
flabel metal4 s 0 7910 200 8840 0 FreeSans 1000 0 0 0 VSSD
port 9 nsew
flabel metal5 s 800 7930 1000 8820 0 FreeSans 1000 0 0 0 VSSD
port 9 nsew
flabel metal4 s 800 7910 1000 8840 0 FreeSans 1000 0 0 0 VSSD
port 9 nsew
flabel metal5 s 0 11260 200 12110 0 FreeSans 1000 0 0 0 VSSIO_Q
port 10 nsew
flabel metal4 s 0 11240 200 12130 0 FreeSans 1000 0 0 0 VSSIO_Q
port 10 nsew
flabel metal5 s 800 11260 1000 12110 0 FreeSans 1000 0 0 0 VSSIO_Q
port 10 nsew
flabel metal4 s 800 11240 1000 12130 0 FreeSans 1000 0 0 0 VSSIO_Q
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 39593
string GDS_END 7104
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_ef_io__disconnect_vdda_slice_5um.gds
string GDS_START 170
<< end >>
