magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 9 -205 12 -202 8 B_P
port 1 nsew
rlabel  s 77 -124 77 -124 8 D_P
port 2 nsew
rlabel  s 76 -124 77 -124 8 D_P
port 2 nsew
rlabel  s 74 -124 81 -124 8 D_P
port 2 nsew
rlabel  s 85 103 97 103 6 G
port 3 nsew
rlabel  s 85 101 85 103 6 G
port 3 nsew
rlabel  s 72 101 85 101 6 G
port 3 nsew
rlabel  s 72 101 73 101 6 G
port 3 nsew
rlabel  s 68 100 73 101 6 G
port 3 nsew
rlabel  s 85 -120 87 -120 8 G_P
port 4 nsew
rlabel  s 85 -122 85 -120 8 G_P
port 4 nsew
rlabel  s 79 -122 85 -122 8 G_P
port 4 nsew
rlabel  s 79 -123 80 -122 8 G_P
port 4 nsew
rlabel  s 76 -123 77 -123 8 G_P
port 4 nsew
rlabel  s 70 -123 80 -123 8 G_P
port 4 nsew
rlabel  s 70 -124 71 -123 8 G_P
port 4 nsew
rlabel  s 67 -124 71 -124 8 G_P
port 4 nsew
rlabel  s 9 9 12 12 6 NWELL
port 5 nsew
rlabel  s 98 100 98 103 6 S
port 6 nsew
rlabel  s 97 100 97 103 6 S
port 6 nsew
rlabel  s 96 100 96 103 6 S
port 6 nsew
rlabel  s 95 100 95 103 6 S
port 6 nsew
rlabel  s 94 100 94 103 6 S
port 6 nsew
rlabel  s 92 100 92 103 6 S
port 6 nsew
rlabel  s 91 100 91 103 6 S
port 6 nsew
rlabel  s 90 100 90 103 6 S
port 6 nsew
rlabel  s 87 100 88 103 6 S
port 6 nsew
rlabel  s 87 100 87 103 6 S
port 6 nsew
rlabel  s 84 100 84 101 6 S
port 6 nsew
rlabel  s 83 100 83 101 6 S
port 6 nsew
rlabel  s 82 100 82 101 6 S
port 6 nsew
rlabel  s 81 100 81 101 6 S
port 6 nsew
rlabel  s 80 100 80 101 6 S
port 6 nsew
rlabel  s 79 100 79 101 6 S
port 6 nsew
rlabel  s 78 100 78 101 6 S
port 6 nsew
rlabel  s 77 100 77 101 6 S
port 6 nsew
rlabel  s 75 100 75 101 6 S
port 6 nsew
rlabel  s 74 100 74 101 6 S
port 6 nsew
rlabel  s 70 100 70 100 6 S
port 6 nsew
rlabel  s 69 100 69 100 6 S
port 6 nsew
rlabel  s 68 99 98 100 6 S
port 6 nsew
rlabel  s 87 -126 87 -120 8 S_P
port 7 nsew
rlabel  s 86 -126 87 -120 8 S_P
port 7 nsew
rlabel  s 83 -126 83 -122 8 S_P
port 7 nsew
rlabel  s 82 -126 82 -122 8 S_P
port 7 nsew
rlabel  s 78 -126 78 -124 8 S_P
port 7 nsew
rlabel  s 77 -126 77 -124 8 S_P
port 7 nsew
rlabel  s 76 -126 76 -124 8 S_P
port 7 nsew
rlabel  s 73 -126 73 -124 8 S_P
port 7 nsew
rlabel  s 72 -126 72 -124 8 S_P
port 7 nsew
rlabel  s 69 -126 69 -125 8 S_P
port 7 nsew
rlabel  s 68 -126 68 -125 8 S_P
port 7 nsew
rlabel  s 67 -126 87 -126 8 S_P
port 7 nsew
rlabel  s 60 91 63 94 6 VGND
port 8 nsew ground default
rlabel  s 89 102 97 103 6 VPWR
port 9 nsew power default
rlabel  s 86 101 86 103 6 VPWR
port 9 nsew power default
rlabel  s 83 100 83 100 6 VPWR
port 9 nsew power default
rlabel  s 82 100 83 100 6 VPWR
port 9 nsew power default
rlabel  s 81 100 82 100 6 VPWR
port 9 nsew power default
rlabel  s 80 100 81 100 6 VPWR
port 9 nsew power default
rlabel  s 78 100 78 100 6 VPWR
port 9 nsew power default
rlabel  s 77 100 78 100 6 VPWR
port 9 nsew power default
rlabel  s 76 100 86 101 6 VPWR
port 9 nsew power default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 -214 1556 198
string LEFview TRUE
<< end >>
