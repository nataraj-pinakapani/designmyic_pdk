magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< pwell >>
rect 10 10 1248 1340
<< mvnmos >>
rect 229 144 1029 1144
<< mvndiff >>
rect 176 1074 229 1144
rect 176 1040 184 1074
rect 218 1040 229 1074
rect 176 1006 229 1040
rect 176 972 184 1006
rect 218 972 229 1006
rect 176 938 229 972
rect 176 904 184 938
rect 218 904 229 938
rect 176 870 229 904
rect 176 836 184 870
rect 218 836 229 870
rect 176 802 229 836
rect 176 768 184 802
rect 218 768 229 802
rect 176 734 229 768
rect 176 700 184 734
rect 218 700 229 734
rect 176 666 229 700
rect 176 632 184 666
rect 218 632 229 666
rect 176 598 229 632
rect 176 564 184 598
rect 218 564 229 598
rect 176 530 229 564
rect 176 496 184 530
rect 218 496 229 530
rect 176 462 229 496
rect 176 428 184 462
rect 218 428 229 462
rect 176 394 229 428
rect 176 360 184 394
rect 218 360 229 394
rect 176 326 229 360
rect 176 292 184 326
rect 218 292 229 326
rect 176 258 229 292
rect 176 224 184 258
rect 218 224 229 258
rect 176 190 229 224
rect 176 156 184 190
rect 218 156 229 190
rect 176 144 229 156
rect 1029 1074 1082 1144
rect 1029 1040 1040 1074
rect 1074 1040 1082 1074
rect 1029 1006 1082 1040
rect 1029 972 1040 1006
rect 1074 972 1082 1006
rect 1029 938 1082 972
rect 1029 904 1040 938
rect 1074 904 1082 938
rect 1029 870 1082 904
rect 1029 836 1040 870
rect 1074 836 1082 870
rect 1029 802 1082 836
rect 1029 768 1040 802
rect 1074 768 1082 802
rect 1029 734 1082 768
rect 1029 700 1040 734
rect 1074 700 1082 734
rect 1029 666 1082 700
rect 1029 632 1040 666
rect 1074 632 1082 666
rect 1029 598 1082 632
rect 1029 564 1040 598
rect 1074 564 1082 598
rect 1029 530 1082 564
rect 1029 496 1040 530
rect 1074 496 1082 530
rect 1029 462 1082 496
rect 1029 428 1040 462
rect 1074 428 1082 462
rect 1029 394 1082 428
rect 1029 360 1040 394
rect 1074 360 1082 394
rect 1029 326 1082 360
rect 1029 292 1040 326
rect 1074 292 1082 326
rect 1029 258 1082 292
rect 1029 224 1040 258
rect 1074 224 1082 258
rect 1029 190 1082 224
rect 1029 156 1040 190
rect 1074 156 1082 190
rect 1029 144 1082 156
<< mvndiffc >>
rect 184 1040 218 1074
rect 184 972 218 1006
rect 184 904 218 938
rect 184 836 218 870
rect 184 768 218 802
rect 184 700 218 734
rect 184 632 218 666
rect 184 564 218 598
rect 184 496 218 530
rect 184 428 218 462
rect 184 360 218 394
rect 184 292 218 326
rect 184 224 218 258
rect 184 156 218 190
rect 1040 1040 1074 1074
rect 1040 972 1074 1006
rect 1040 904 1074 938
rect 1040 836 1074 870
rect 1040 768 1074 802
rect 1040 700 1074 734
rect 1040 632 1074 666
rect 1040 564 1074 598
rect 1040 496 1074 530
rect 1040 428 1074 462
rect 1040 360 1074 394
rect 1040 292 1074 326
rect 1040 224 1074 258
rect 1040 156 1074 190
<< mvpsubdiff >>
rect 36 1246 70 1314
rect 104 1280 138 1314
rect 172 1280 206 1314
rect 240 1280 274 1314
rect 308 1280 342 1314
rect 376 1280 410 1314
rect 444 1280 478 1314
rect 512 1280 546 1314
rect 580 1280 614 1314
rect 648 1280 682 1314
rect 716 1280 750 1314
rect 784 1280 818 1314
rect 852 1280 886 1314
rect 920 1280 954 1314
rect 988 1280 1022 1314
rect 1056 1280 1090 1314
rect 1124 1280 1222 1314
rect 1188 1246 1222 1280
rect 36 1178 70 1212
rect 1188 1178 1222 1212
rect 36 1110 70 1144
rect 36 1042 70 1076
rect 36 974 70 1008
rect 36 906 70 940
rect 36 838 70 872
rect 36 770 70 804
rect 36 702 70 736
rect 36 634 70 668
rect 36 566 70 600
rect 36 498 70 532
rect 36 430 70 464
rect 36 362 70 396
rect 36 294 70 328
rect 36 226 70 260
rect 36 158 70 192
rect 1188 1110 1222 1144
rect 1188 1042 1222 1076
rect 1188 974 1222 1008
rect 1188 906 1222 940
rect 1188 838 1222 872
rect 1188 770 1222 804
rect 1188 702 1222 736
rect 1188 634 1222 668
rect 1188 566 1222 600
rect 1188 498 1222 532
rect 1188 430 1222 464
rect 1188 362 1222 396
rect 1188 294 1222 328
rect 1188 226 1222 260
rect 1188 158 1222 192
rect 36 36 70 124
rect 1188 70 1222 124
rect 104 36 138 70
rect 172 36 206 70
rect 240 36 274 70
rect 308 36 342 70
rect 376 36 410 70
rect 444 36 478 70
rect 512 36 546 70
rect 580 36 614 70
rect 648 36 682 70
rect 716 36 750 70
rect 784 36 818 70
rect 852 36 886 70
rect 920 36 954 70
rect 988 36 1022 70
rect 1056 36 1090 70
rect 1124 36 1222 70
<< mvpsubdiffcont >>
rect 70 1280 104 1314
rect 138 1280 172 1314
rect 206 1280 240 1314
rect 274 1280 308 1314
rect 342 1280 376 1314
rect 410 1280 444 1314
rect 478 1280 512 1314
rect 546 1280 580 1314
rect 614 1280 648 1314
rect 682 1280 716 1314
rect 750 1280 784 1314
rect 818 1280 852 1314
rect 886 1280 920 1314
rect 954 1280 988 1314
rect 1022 1280 1056 1314
rect 1090 1280 1124 1314
rect 36 1212 70 1246
rect 36 1144 70 1178
rect 1188 1212 1222 1246
rect 1188 1144 1222 1178
rect 36 1076 70 1110
rect 36 1008 70 1042
rect 36 940 70 974
rect 36 872 70 906
rect 36 804 70 838
rect 36 736 70 770
rect 36 668 70 702
rect 36 600 70 634
rect 36 532 70 566
rect 36 464 70 498
rect 36 396 70 430
rect 36 328 70 362
rect 36 260 70 294
rect 36 192 70 226
rect 36 124 70 158
rect 1188 1076 1222 1110
rect 1188 1008 1222 1042
rect 1188 940 1222 974
rect 1188 872 1222 906
rect 1188 804 1222 838
rect 1188 736 1222 770
rect 1188 668 1222 702
rect 1188 600 1222 634
rect 1188 532 1222 566
rect 1188 464 1222 498
rect 1188 396 1222 430
rect 1188 328 1222 362
rect 1188 260 1222 294
rect 1188 192 1222 226
rect 1188 124 1222 158
rect 70 36 104 70
rect 138 36 172 70
rect 206 36 240 70
rect 274 36 308 70
rect 342 36 376 70
rect 410 36 444 70
rect 478 36 512 70
rect 546 36 580 70
rect 614 36 648 70
rect 682 36 716 70
rect 750 36 784 70
rect 818 36 852 70
rect 886 36 920 70
rect 954 36 988 70
rect 1022 36 1056 70
rect 1090 36 1124 70
<< poly >>
rect 229 1220 1029 1236
rect 229 1186 249 1220
rect 283 1186 317 1220
rect 351 1186 385 1220
rect 419 1186 453 1220
rect 487 1186 521 1220
rect 555 1186 589 1220
rect 623 1186 657 1220
rect 691 1186 725 1220
rect 759 1186 793 1220
rect 827 1186 861 1220
rect 895 1186 929 1220
rect 963 1186 1029 1220
rect 229 1144 1029 1186
rect 229 118 1029 144
<< polycont >>
rect 249 1186 283 1220
rect 317 1186 351 1220
rect 385 1186 419 1220
rect 453 1186 487 1220
rect 521 1186 555 1220
rect 589 1186 623 1220
rect 657 1186 691 1220
rect 725 1186 759 1220
rect 793 1186 827 1220
rect 861 1186 895 1220
rect 929 1186 963 1220
<< locali >>
rect 70 1314 1188 1320
rect 36 1280 70 1314
rect 116 1280 138 1314
rect 188 1280 206 1314
rect 260 1280 274 1314
rect 332 1280 342 1314
rect 404 1280 410 1314
rect 476 1280 478 1314
rect 512 1280 514 1314
rect 580 1280 586 1314
rect 648 1280 658 1314
rect 716 1280 730 1314
rect 784 1280 802 1314
rect 852 1280 874 1314
rect 920 1280 946 1314
rect 988 1280 1018 1314
rect 1056 1280 1090 1314
rect 1124 1280 1222 1314
rect 36 1274 1222 1280
rect 36 1246 70 1274
rect 1188 1246 1222 1274
rect 36 1178 70 1212
rect 229 1220 1029 1226
rect 229 1186 241 1220
rect 283 1186 313 1220
rect 351 1186 385 1220
rect 419 1186 453 1220
rect 491 1186 521 1220
rect 563 1186 589 1220
rect 635 1186 657 1220
rect 707 1186 725 1220
rect 779 1186 793 1220
rect 851 1186 861 1220
rect 923 1186 929 1220
rect 995 1186 1029 1220
rect 229 1180 1029 1186
rect 36 1110 70 1144
rect 1188 1178 1222 1212
rect 1188 1110 1222 1144
rect 36 1042 70 1076
rect 36 974 70 1008
rect 36 906 70 940
rect 30 872 36 877
rect 184 1074 218 1090
rect 184 1006 218 1040
rect 184 938 218 972
rect 184 877 218 904
rect 1040 1074 1074 1090
rect 1040 1006 1074 1040
rect 1040 938 1074 972
rect 1040 877 1074 904
rect 1188 1042 1222 1076
rect 1188 974 1222 1008
rect 1188 906 1222 940
rect 70 872 76 877
rect 30 865 76 872
rect 30 804 36 865
rect 70 804 76 865
rect 30 793 76 804
rect 30 736 36 793
rect 70 736 76 793
rect 30 721 76 736
rect 30 668 36 721
rect 70 668 76 721
rect 30 649 76 668
rect 30 600 36 649
rect 70 600 76 649
rect 30 577 76 600
rect 30 532 36 577
rect 70 532 76 577
rect 30 505 76 532
rect 30 464 36 505
rect 70 464 76 505
rect 30 433 76 464
rect 30 396 36 433
rect 70 396 76 433
rect 30 362 76 396
rect 30 327 36 362
rect 70 327 76 362
rect 30 294 76 327
rect 30 255 36 294
rect 70 255 76 294
rect 176 870 222 877
rect 176 865 184 870
rect 176 831 182 865
rect 218 836 222 870
rect 216 831 222 836
rect 176 802 222 831
rect 176 793 184 802
rect 176 759 182 793
rect 218 768 222 802
rect 216 759 222 768
rect 176 734 222 759
rect 176 721 184 734
rect 176 687 182 721
rect 218 700 222 734
rect 216 687 222 700
rect 176 666 222 687
rect 176 649 184 666
rect 176 615 182 649
rect 218 632 222 666
rect 216 615 222 632
rect 176 598 222 615
rect 176 577 184 598
rect 176 543 182 577
rect 218 564 222 598
rect 216 543 222 564
rect 176 530 222 543
rect 176 505 184 530
rect 176 471 182 505
rect 218 496 222 530
rect 216 471 222 496
rect 176 462 222 471
rect 176 433 184 462
rect 176 399 182 433
rect 218 428 222 462
rect 216 399 222 428
rect 176 394 222 399
rect 176 361 184 394
rect 176 327 182 361
rect 218 360 222 394
rect 216 327 222 360
rect 176 326 222 327
rect 176 292 184 326
rect 218 292 222 326
rect 176 287 222 292
rect 1035 870 1081 877
rect 1035 836 1040 870
rect 1074 865 1081 870
rect 1035 831 1041 836
rect 1075 831 1081 865
rect 1035 802 1081 831
rect 1035 768 1040 802
rect 1074 793 1081 802
rect 1035 759 1041 768
rect 1075 759 1081 793
rect 1035 734 1081 759
rect 1035 700 1040 734
rect 1074 721 1081 734
rect 1035 687 1041 700
rect 1075 687 1081 721
rect 1035 666 1081 687
rect 1035 632 1040 666
rect 1074 649 1081 666
rect 1035 615 1041 632
rect 1075 615 1081 649
rect 1035 598 1081 615
rect 1035 564 1040 598
rect 1074 577 1081 598
rect 1035 543 1041 564
rect 1075 543 1081 577
rect 1035 530 1081 543
rect 1035 496 1040 530
rect 1074 505 1081 530
rect 1035 471 1041 496
rect 1075 471 1081 505
rect 1035 462 1081 471
rect 1035 428 1040 462
rect 1074 433 1081 462
rect 1035 399 1041 428
rect 1075 399 1081 433
rect 1035 394 1081 399
rect 1035 360 1040 394
rect 1074 361 1081 394
rect 1035 327 1041 360
rect 1075 327 1081 361
rect 1035 326 1081 327
rect 1035 292 1040 326
rect 1074 292 1081 326
rect 1035 287 1081 292
rect 1182 872 1188 877
rect 1222 872 1228 877
rect 1182 865 1228 872
rect 1182 804 1188 865
rect 1222 804 1228 865
rect 1182 793 1228 804
rect 1182 736 1188 793
rect 1222 736 1228 793
rect 1182 721 1228 736
rect 1182 668 1188 721
rect 1222 668 1228 721
rect 1182 649 1228 668
rect 1182 600 1188 649
rect 1222 600 1228 649
rect 1182 577 1228 600
rect 1182 532 1188 577
rect 1222 532 1228 577
rect 1182 505 1228 532
rect 1182 464 1188 505
rect 1222 464 1228 505
rect 1182 433 1228 464
rect 1182 396 1188 433
rect 1222 396 1228 433
rect 1182 362 1228 396
rect 1182 327 1188 362
rect 1222 327 1228 362
rect 1182 294 1228 327
rect 30 226 76 255
rect 30 183 36 226
rect 70 183 76 226
rect 30 158 76 183
rect 30 111 36 158
rect 70 111 76 158
rect 184 258 218 287
rect 184 190 218 224
rect 184 140 218 156
rect 1040 258 1074 287
rect 1040 190 1074 224
rect 1040 140 1074 156
rect 1182 255 1188 294
rect 1222 255 1228 294
rect 1182 226 1228 255
rect 1182 183 1188 226
rect 1222 183 1228 226
rect 1182 158 1228 183
rect 30 76 76 111
rect 1182 111 1188 158
rect 1222 111 1228 158
rect 1182 76 1228 111
rect 30 70 1228 76
rect 30 36 70 70
rect 116 36 138 70
rect 188 36 206 70
rect 260 36 274 70
rect 332 36 342 70
rect 404 36 410 70
rect 476 36 478 70
rect 512 36 514 70
rect 580 36 586 70
rect 648 36 658 70
rect 716 36 730 70
rect 784 36 802 70
rect 852 36 874 70
rect 920 36 946 70
rect 988 36 1018 70
rect 1056 36 1090 70
rect 1124 36 1228 70
rect 30 30 1228 36
<< viali >>
rect 82 1280 104 1314
rect 104 1280 116 1314
rect 154 1280 172 1314
rect 172 1280 188 1314
rect 226 1280 240 1314
rect 240 1280 260 1314
rect 298 1280 308 1314
rect 308 1280 332 1314
rect 370 1280 376 1314
rect 376 1280 404 1314
rect 442 1280 444 1314
rect 444 1280 476 1314
rect 514 1280 546 1314
rect 546 1280 548 1314
rect 586 1280 614 1314
rect 614 1280 620 1314
rect 658 1280 682 1314
rect 682 1280 692 1314
rect 730 1280 750 1314
rect 750 1280 764 1314
rect 802 1280 818 1314
rect 818 1280 836 1314
rect 874 1280 886 1314
rect 886 1280 908 1314
rect 946 1280 954 1314
rect 954 1280 980 1314
rect 1018 1280 1022 1314
rect 1022 1280 1052 1314
rect 1090 1280 1124 1314
rect 241 1186 249 1220
rect 249 1186 275 1220
rect 313 1186 317 1220
rect 317 1186 347 1220
rect 385 1186 419 1220
rect 457 1186 487 1220
rect 487 1186 491 1220
rect 529 1186 555 1220
rect 555 1186 563 1220
rect 601 1186 623 1220
rect 623 1186 635 1220
rect 673 1186 691 1220
rect 691 1186 707 1220
rect 745 1186 759 1220
rect 759 1186 779 1220
rect 817 1186 827 1220
rect 827 1186 851 1220
rect 889 1186 895 1220
rect 895 1186 923 1220
rect 961 1186 963 1220
rect 963 1186 995 1220
rect 36 838 70 865
rect 36 831 70 838
rect 36 770 70 793
rect 36 759 70 770
rect 36 702 70 721
rect 36 687 70 702
rect 36 634 70 649
rect 36 615 70 634
rect 36 566 70 577
rect 36 543 70 566
rect 36 498 70 505
rect 36 471 70 498
rect 36 430 70 433
rect 36 399 70 430
rect 36 328 70 361
rect 36 327 70 328
rect 36 260 70 289
rect 36 255 70 260
rect 182 836 184 865
rect 184 836 216 865
rect 182 831 216 836
rect 182 768 184 793
rect 184 768 216 793
rect 182 759 216 768
rect 182 700 184 721
rect 184 700 216 721
rect 182 687 216 700
rect 182 632 184 649
rect 184 632 216 649
rect 182 615 216 632
rect 182 564 184 577
rect 184 564 216 577
rect 182 543 216 564
rect 182 496 184 505
rect 184 496 216 505
rect 182 471 216 496
rect 182 428 184 433
rect 184 428 216 433
rect 182 399 216 428
rect 182 360 184 361
rect 184 360 216 361
rect 182 327 216 360
rect 1041 836 1074 865
rect 1074 836 1075 865
rect 1041 831 1075 836
rect 1041 768 1074 793
rect 1074 768 1075 793
rect 1041 759 1075 768
rect 1041 700 1074 721
rect 1074 700 1075 721
rect 1041 687 1075 700
rect 1041 632 1074 649
rect 1074 632 1075 649
rect 1041 615 1075 632
rect 1041 564 1074 577
rect 1074 564 1075 577
rect 1041 543 1075 564
rect 1041 496 1074 505
rect 1074 496 1075 505
rect 1041 471 1075 496
rect 1041 428 1074 433
rect 1074 428 1075 433
rect 1041 399 1075 428
rect 1041 360 1074 361
rect 1074 360 1075 361
rect 1041 327 1075 360
rect 1188 838 1222 865
rect 1188 831 1222 838
rect 1188 770 1222 793
rect 1188 759 1222 770
rect 1188 702 1222 721
rect 1188 687 1222 702
rect 1188 634 1222 649
rect 1188 615 1222 634
rect 1188 566 1222 577
rect 1188 543 1222 566
rect 1188 498 1222 505
rect 1188 471 1222 498
rect 1188 430 1222 433
rect 1188 399 1222 430
rect 1188 328 1222 361
rect 1188 327 1222 328
rect 36 192 70 217
rect 36 183 70 192
rect 36 124 70 145
rect 36 111 70 124
rect 1188 260 1222 289
rect 1188 255 1222 260
rect 1188 192 1222 217
rect 1188 183 1222 192
rect 1188 124 1222 145
rect 1188 111 1222 124
rect 82 36 104 70
rect 104 36 116 70
rect 154 36 172 70
rect 172 36 188 70
rect 226 36 240 70
rect 240 36 260 70
rect 298 36 308 70
rect 308 36 332 70
rect 370 36 376 70
rect 376 36 404 70
rect 442 36 444 70
rect 444 36 476 70
rect 514 36 546 70
rect 546 36 548 70
rect 586 36 614 70
rect 614 36 620 70
rect 658 36 682 70
rect 682 36 692 70
rect 730 36 750 70
rect 750 36 764 70
rect 802 36 818 70
rect 818 36 836 70
rect 874 36 886 70
rect 886 36 908 70
rect 946 36 954 70
rect 954 36 980 70
rect 1018 36 1022 70
rect 1022 36 1052 70
rect 1090 36 1124 70
<< metal1 >>
rect 36 1314 1222 1320
rect 36 1280 82 1314
rect 116 1280 154 1314
rect 188 1280 226 1314
rect 260 1280 298 1314
rect 332 1280 370 1314
rect 404 1280 442 1314
rect 476 1280 514 1314
rect 548 1280 586 1314
rect 620 1280 658 1314
rect 692 1280 730 1314
rect 764 1280 802 1314
rect 836 1280 874 1314
rect 908 1280 946 1314
rect 980 1280 1018 1314
rect 1052 1280 1090 1314
rect 1124 1280 1222 1314
rect 36 1274 1222 1280
rect 28 1220 1230 1229
rect 28 1186 241 1220
rect 275 1186 313 1220
rect 347 1186 385 1220
rect 419 1186 457 1220
rect 491 1186 529 1220
rect 563 1186 601 1220
rect 635 1186 673 1220
rect 707 1186 745 1220
rect 779 1186 817 1220
rect 851 1186 889 1220
rect 923 1186 961 1220
rect 995 1186 1230 1220
rect 28 1177 1230 1186
rect 30 865 1228 877
rect 30 831 36 865
rect 70 831 182 865
rect 216 831 1041 865
rect 1075 831 1188 865
rect 1222 831 1228 865
rect 30 793 1228 831
rect 30 759 36 793
rect 70 759 182 793
rect 216 759 1041 793
rect 1075 759 1188 793
rect 1222 759 1228 793
rect 30 721 1228 759
rect 30 687 36 721
rect 70 687 182 721
rect 216 687 1041 721
rect 1075 687 1188 721
rect 1222 687 1228 721
rect 30 649 1228 687
rect 30 615 36 649
rect 70 615 182 649
rect 216 615 1041 649
rect 1075 615 1188 649
rect 1222 615 1228 649
rect 30 577 1228 615
rect 30 543 36 577
rect 70 543 182 577
rect 216 543 1041 577
rect 1075 543 1188 577
rect 1222 543 1228 577
rect 30 505 1228 543
rect 30 471 36 505
rect 70 471 182 505
rect 216 471 1041 505
rect 1075 471 1188 505
rect 1222 471 1228 505
rect 30 433 1228 471
rect 30 399 36 433
rect 70 399 182 433
rect 216 399 1041 433
rect 1075 399 1188 433
rect 1222 399 1228 433
rect 30 361 1228 399
rect 30 327 36 361
rect 70 327 182 361
rect 216 327 1041 361
rect 1075 327 1188 361
rect 1222 327 1228 361
rect 30 289 1228 327
rect 30 255 36 289
rect 70 287 1188 289
rect 70 255 78 287
tri 78 255 110 287 nw
tri 1148 255 1180 287 ne
rect 1180 255 1188 287
rect 1222 255 1228 289
rect 30 217 76 255
tri 76 253 78 255 nw
tri 1180 253 1182 255 ne
rect 30 183 36 217
rect 70 183 76 217
rect 30 145 76 183
rect 30 111 36 145
rect 70 111 76 145
rect 30 76 76 111
rect 1182 217 1228 255
rect 1182 183 1188 217
rect 1222 183 1228 217
rect 1182 145 1228 183
rect 1182 111 1188 145
rect 1222 111 1228 145
tri 76 76 110 110 sw
tri 1148 76 1182 110 se
rect 1182 76 1228 111
rect 30 70 1228 76
rect 30 36 82 70
rect 116 36 154 70
rect 188 36 226 70
rect 260 36 298 70
rect 332 36 370 70
rect 404 36 442 70
rect 476 36 514 70
rect 548 36 586 70
rect 620 36 658 70
rect 692 36 730 70
rect 764 36 802 70
rect 836 36 874 70
rect 908 36 946 70
rect 980 36 1018 70
rect 1052 36 1090 70
rect 1124 36 1228 70
rect 30 30 1228 36
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808664  sky130_fd_pr__model__nfet_highvoltage__example_55959141808664_0
timestamp 1663361622
transform 1 0 229 0 1 144
box -1 0 801 1
<< properties >>
string GDS_END 11803768
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 11790910
<< end >>
