magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 0 0 776 806
<< pmos >>
rect 204 102 254 704
rect 310 102 360 704
rect 416 102 466 704
rect 522 102 572 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 254 692 310 704
rect 254 658 265 692
rect 299 658 310 692
rect 254 624 310 658
rect 254 590 265 624
rect 299 590 310 624
rect 254 556 310 590
rect 254 522 265 556
rect 299 522 310 556
rect 254 488 310 522
rect 254 454 265 488
rect 299 454 310 488
rect 254 420 310 454
rect 254 386 265 420
rect 299 386 310 420
rect 254 352 310 386
rect 254 318 265 352
rect 299 318 310 352
rect 254 284 310 318
rect 254 250 265 284
rect 299 250 310 284
rect 254 216 310 250
rect 254 182 265 216
rect 299 182 310 216
rect 254 148 310 182
rect 254 114 265 148
rect 299 114 310 148
rect 254 102 310 114
rect 360 692 416 704
rect 360 658 371 692
rect 405 658 416 692
rect 360 624 416 658
rect 360 590 371 624
rect 405 590 416 624
rect 360 556 416 590
rect 360 522 371 556
rect 405 522 416 556
rect 360 488 416 522
rect 360 454 371 488
rect 405 454 416 488
rect 360 420 416 454
rect 360 386 371 420
rect 405 386 416 420
rect 360 352 416 386
rect 360 318 371 352
rect 405 318 416 352
rect 360 284 416 318
rect 360 250 371 284
rect 405 250 416 284
rect 360 216 416 250
rect 360 182 371 216
rect 405 182 416 216
rect 360 148 416 182
rect 360 114 371 148
rect 405 114 416 148
rect 360 102 416 114
rect 466 692 522 704
rect 466 658 477 692
rect 511 658 522 692
rect 466 624 522 658
rect 466 590 477 624
rect 511 590 522 624
rect 466 556 522 590
rect 466 522 477 556
rect 511 522 522 556
rect 466 488 522 522
rect 466 454 477 488
rect 511 454 522 488
rect 466 420 522 454
rect 466 386 477 420
rect 511 386 522 420
rect 466 352 522 386
rect 466 318 477 352
rect 511 318 522 352
rect 466 284 522 318
rect 466 250 477 284
rect 511 250 522 284
rect 466 216 522 250
rect 466 182 477 216
rect 511 182 522 216
rect 466 148 522 182
rect 466 114 477 148
rect 511 114 522 148
rect 466 102 522 114
rect 572 692 628 704
rect 572 658 583 692
rect 617 658 628 692
rect 572 624 628 658
rect 572 590 583 624
rect 617 590 628 624
rect 572 556 628 590
rect 572 522 583 556
rect 617 522 628 556
rect 572 488 628 522
rect 572 454 583 488
rect 617 454 628 488
rect 572 420 628 454
rect 572 386 583 420
rect 617 386 628 420
rect 572 352 628 386
rect 572 318 583 352
rect 617 318 628 352
rect 572 284 628 318
rect 572 250 583 284
rect 617 250 628 284
rect 572 216 628 250
rect 572 182 583 216
rect 617 182 628 216
rect 572 148 628 182
rect 572 114 583 148
rect 617 114 628 148
rect 572 102 628 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 265 658 299 692
rect 265 590 299 624
rect 265 522 299 556
rect 265 454 299 488
rect 265 386 299 420
rect 265 318 299 352
rect 265 250 299 284
rect 265 182 299 216
rect 265 114 299 148
rect 371 658 405 692
rect 371 590 405 624
rect 371 522 405 556
rect 371 454 405 488
rect 371 386 405 420
rect 371 318 405 352
rect 371 250 405 284
rect 371 182 405 216
rect 371 114 405 148
rect 477 658 511 692
rect 477 590 511 624
rect 477 522 511 556
rect 477 454 511 488
rect 477 386 511 420
rect 477 318 511 352
rect 477 250 511 284
rect 477 182 511 216
rect 477 114 511 148
rect 583 658 617 692
rect 583 590 617 624
rect 583 522 617 556
rect 583 454 617 488
rect 583 386 617 420
rect 583 318 617 352
rect 583 250 617 284
rect 583 182 617 216
rect 583 114 617 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 682 658 740 704
rect 682 624 694 658
rect 728 624 740 658
rect 682 590 740 624
rect 682 556 694 590
rect 728 556 740 590
rect 682 522 740 556
rect 682 488 694 522
rect 728 488 740 522
rect 682 454 740 488
rect 682 420 694 454
rect 728 420 740 454
rect 682 386 740 420
rect 682 352 694 386
rect 728 352 740 386
rect 682 318 740 352
rect 682 284 694 318
rect 728 284 740 318
rect 682 250 740 284
rect 682 216 694 250
rect 728 216 740 250
rect 682 182 740 216
rect 682 148 694 182
rect 728 148 740 182
rect 682 102 740 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 694 624 728 658
rect 694 556 728 590
rect 694 488 728 522
rect 694 420 728 454
rect 694 352 728 386
rect 694 284 728 318
rect 694 216 728 250
rect 694 148 728 182
<< poly >>
rect 185 786 591 806
rect 185 752 201 786
rect 235 752 269 786
rect 303 752 337 786
rect 371 752 405 786
rect 439 752 473 786
rect 507 752 541 786
rect 575 752 591 786
rect 185 736 591 752
rect 204 704 254 736
rect 310 704 360 736
rect 416 704 466 736
rect 522 704 572 736
rect 204 70 254 102
rect 310 70 360 102
rect 416 70 466 102
rect 522 70 572 102
rect 185 54 591 70
rect 185 20 201 54
rect 235 20 269 54
rect 303 20 337 54
rect 371 20 405 54
rect 439 20 473 54
rect 507 20 541 54
rect 575 20 591 54
rect 185 0 591 20
<< polycont >>
rect 201 752 235 786
rect 269 752 303 786
rect 337 752 371 786
rect 405 752 439 786
rect 473 752 507 786
rect 541 752 575 786
rect 201 20 235 54
rect 269 20 303 54
rect 337 20 371 54
rect 405 20 439 54
rect 473 20 507 54
rect 541 20 575 54
<< locali >>
rect 185 752 192 786
rect 235 752 264 786
rect 303 752 336 786
rect 371 752 405 786
rect 442 752 473 786
rect 514 752 541 786
rect 586 752 591 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 265 692 299 708
rect 265 624 299 638
rect 265 556 299 566
rect 265 488 299 494
rect 265 420 299 422
rect 265 384 299 386
rect 265 312 299 318
rect 265 240 299 250
rect 265 168 299 182
rect 265 98 299 114
rect 371 692 405 708
rect 371 624 405 638
rect 371 556 405 566
rect 371 488 405 494
rect 371 420 405 422
rect 371 384 405 386
rect 371 312 405 318
rect 371 240 405 250
rect 371 168 405 182
rect 371 98 405 114
rect 477 692 511 708
rect 477 624 511 638
rect 477 556 511 566
rect 477 488 511 494
rect 477 420 511 422
rect 477 384 511 386
rect 477 312 511 318
rect 477 240 511 250
rect 477 168 511 182
rect 477 98 511 114
rect 583 692 617 708
rect 583 624 617 638
rect 583 556 617 566
rect 583 488 617 494
rect 583 420 617 422
rect 583 384 617 386
rect 583 312 617 318
rect 583 240 617 250
rect 583 168 617 182
rect 694 672 728 674
rect 694 600 728 624
rect 694 528 728 556
rect 694 456 728 488
rect 694 386 728 420
rect 694 318 728 350
rect 694 250 728 278
rect 694 182 728 206
rect 694 132 728 134
rect 583 98 617 114
rect 185 20 192 54
rect 235 20 264 54
rect 303 20 336 54
rect 371 20 405 54
rect 442 20 473 54
rect 514 20 541 54
rect 586 20 591 54
<< viali >>
rect 192 752 201 786
rect 201 752 226 786
rect 264 752 269 786
rect 269 752 298 786
rect 336 752 337 786
rect 337 752 370 786
rect 408 752 439 786
rect 439 752 442 786
rect 480 752 507 786
rect 507 752 514 786
rect 552 752 575 786
rect 575 752 586 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 265 658 299 672
rect 265 638 299 658
rect 265 590 299 600
rect 265 566 299 590
rect 265 522 299 528
rect 265 494 299 522
rect 265 454 299 456
rect 265 422 299 454
rect 265 352 299 384
rect 265 350 299 352
rect 265 284 299 312
rect 265 278 299 284
rect 265 216 299 240
rect 265 206 299 216
rect 265 148 299 168
rect 265 134 299 148
rect 371 658 405 672
rect 371 638 405 658
rect 371 590 405 600
rect 371 566 405 590
rect 371 522 405 528
rect 371 494 405 522
rect 371 454 405 456
rect 371 422 405 454
rect 371 352 405 384
rect 371 350 405 352
rect 371 284 405 312
rect 371 278 405 284
rect 371 216 405 240
rect 371 206 405 216
rect 371 148 405 168
rect 371 134 405 148
rect 477 658 511 672
rect 477 638 511 658
rect 477 590 511 600
rect 477 566 511 590
rect 477 522 511 528
rect 477 494 511 522
rect 477 454 511 456
rect 477 422 511 454
rect 477 352 511 384
rect 477 350 511 352
rect 477 284 511 312
rect 477 278 511 284
rect 477 216 511 240
rect 477 206 511 216
rect 477 148 511 168
rect 477 134 511 148
rect 583 658 617 672
rect 583 638 617 658
rect 583 590 617 600
rect 583 566 617 590
rect 583 522 617 528
rect 583 494 617 522
rect 583 454 617 456
rect 583 422 617 454
rect 583 352 617 384
rect 583 350 617 352
rect 583 284 617 312
rect 583 278 617 284
rect 583 216 617 240
rect 583 206 617 216
rect 583 148 617 168
rect 583 134 617 148
rect 694 658 728 672
rect 694 638 728 658
rect 694 590 728 600
rect 694 566 728 590
rect 694 522 728 528
rect 694 494 728 522
rect 694 454 728 456
rect 694 422 728 454
rect 694 352 728 384
rect 694 350 728 352
rect 694 284 728 312
rect 694 278 728 284
rect 694 216 728 240
rect 694 206 728 216
rect 694 148 728 168
rect 694 134 728 148
rect 192 20 201 54
rect 201 20 226 54
rect 264 20 269 54
rect 269 20 298 54
rect 336 20 337 54
rect 337 20 370 54
rect 408 20 439 54
rect 439 20 442 54
rect 480 20 507 54
rect 507 20 514 54
rect 552 20 575 54
rect 575 20 586 54
<< metal1 >>
rect 180 786 598 806
rect 180 752 192 786
rect 226 752 264 786
rect 298 752 336 786
rect 370 752 408 786
rect 442 752 480 786
rect 514 752 552 786
rect 586 752 598 786
rect 180 740 598 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 256 678 308 684
rect 256 614 308 626
rect 256 550 308 562
rect 256 494 265 498
rect 299 494 308 498
rect 256 486 308 494
rect 256 422 265 434
rect 299 422 308 434
rect 256 384 308 422
rect 256 350 265 384
rect 299 350 308 384
rect 256 312 308 350
rect 256 278 265 312
rect 299 278 308 312
rect 256 240 308 278
rect 256 206 265 240
rect 299 206 308 240
rect 256 168 308 206
rect 256 134 265 168
rect 299 134 308 168
rect 256 122 308 134
rect 362 672 414 684
rect 362 638 371 672
rect 405 638 414 672
rect 362 600 414 638
rect 362 566 371 600
rect 405 566 414 600
rect 362 528 414 566
rect 362 494 371 528
rect 405 494 414 528
rect 362 456 414 494
rect 362 422 371 456
rect 405 422 414 456
rect 362 384 414 422
rect 362 372 371 384
rect 405 372 414 384
rect 362 312 414 320
rect 362 308 371 312
rect 405 308 414 312
rect 362 244 414 256
rect 362 180 414 192
rect 362 122 414 128
rect 468 678 520 684
rect 468 614 520 626
rect 468 550 520 562
rect 468 494 477 498
rect 511 494 520 498
rect 468 486 520 494
rect 468 422 477 434
rect 511 422 520 434
rect 468 384 520 422
rect 468 350 477 384
rect 511 350 520 384
rect 468 312 520 350
rect 468 278 477 312
rect 511 278 520 312
rect 468 240 520 278
rect 468 206 477 240
rect 511 206 520 240
rect 468 168 520 206
rect 468 134 477 168
rect 511 134 520 168
rect 468 122 520 134
rect 574 672 626 684
rect 574 638 583 672
rect 617 638 626 672
rect 574 600 626 638
rect 574 566 583 600
rect 617 566 626 600
rect 574 528 626 566
rect 574 494 583 528
rect 617 494 626 528
rect 574 456 626 494
rect 574 422 583 456
rect 617 422 626 456
rect 574 384 626 422
rect 574 372 583 384
rect 617 372 626 384
rect 574 312 626 320
rect 574 308 583 312
rect 617 308 626 312
rect 574 244 626 256
rect 574 180 626 192
rect 574 122 626 128
rect 682 672 740 684
rect 682 638 694 672
rect 728 638 740 672
rect 682 600 740 638
rect 682 566 694 600
rect 728 566 740 600
rect 682 528 740 566
rect 682 494 694 528
rect 728 494 740 528
rect 682 456 740 494
rect 682 422 694 456
rect 728 422 740 456
rect 682 384 740 422
rect 682 350 694 384
rect 728 350 740 384
rect 682 312 740 350
rect 682 278 694 312
rect 728 278 740 312
rect 682 240 740 278
rect 682 206 694 240
rect 728 206 740 240
rect 682 168 740 206
rect 682 134 694 168
rect 728 134 740 168
rect 682 122 740 134
rect 180 54 598 66
rect 180 20 192 54
rect 226 20 264 54
rect 298 20 336 54
rect 370 20 408 54
rect 442 20 480 54
rect 514 20 552 54
rect 586 20 598 54
rect 180 0 598 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 256 672 308 678
rect 256 638 265 672
rect 265 638 299 672
rect 299 638 308 672
rect 256 626 308 638
rect 256 600 308 614
rect 256 566 265 600
rect 265 566 299 600
rect 299 566 308 600
rect 256 562 308 566
rect 256 528 308 550
rect 256 498 265 528
rect 265 498 299 528
rect 299 498 308 528
rect 256 456 308 486
rect 256 434 265 456
rect 265 434 299 456
rect 299 434 308 456
rect 362 350 371 372
rect 371 350 405 372
rect 405 350 414 372
rect 362 320 414 350
rect 362 278 371 308
rect 371 278 405 308
rect 405 278 414 308
rect 362 256 414 278
rect 362 240 414 244
rect 362 206 371 240
rect 371 206 405 240
rect 405 206 414 240
rect 362 192 414 206
rect 362 168 414 180
rect 362 134 371 168
rect 371 134 405 168
rect 405 134 414 168
rect 362 128 414 134
rect 468 672 520 678
rect 468 638 477 672
rect 477 638 511 672
rect 511 638 520 672
rect 468 626 520 638
rect 468 600 520 614
rect 468 566 477 600
rect 477 566 511 600
rect 511 566 520 600
rect 468 562 520 566
rect 468 528 520 550
rect 468 498 477 528
rect 477 498 511 528
rect 511 498 520 528
rect 468 456 520 486
rect 468 434 477 456
rect 477 434 511 456
rect 511 434 520 456
rect 574 350 583 372
rect 583 350 617 372
rect 617 350 626 372
rect 574 320 626 350
rect 574 278 583 308
rect 583 278 617 308
rect 617 278 626 308
rect 574 256 626 278
rect 574 240 626 244
rect 574 206 583 240
rect 583 206 617 240
rect 617 206 626 240
rect 574 192 626 206
rect 574 168 626 180
rect 574 134 583 168
rect 583 134 617 168
rect 617 134 626 168
rect 574 128 626 134
<< metal2 >>
rect 10 678 766 684
rect 10 626 256 678
rect 308 626 468 678
rect 520 626 766 678
rect 10 614 766 626
rect 10 562 256 614
rect 308 562 468 614
rect 520 562 766 614
rect 10 550 766 562
rect 10 498 256 550
rect 308 498 468 550
rect 520 498 766 550
rect 10 486 766 498
rect 10 434 256 486
rect 308 434 468 486
rect 520 434 766 486
rect 10 428 766 434
rect 10 372 766 378
rect 10 320 150 372
rect 202 320 362 372
rect 414 320 574 372
rect 626 320 766 372
rect 10 308 766 320
rect 10 256 150 308
rect 202 256 362 308
rect 414 256 574 308
rect 626 256 766 308
rect 10 244 766 256
rect 10 192 150 244
rect 202 192 362 244
rect 414 192 574 244
rect 626 192 766 244
rect 10 180 766 192
rect 10 128 150 180
rect 202 128 362 180
rect 414 128 574 180
rect 626 128 766 180
rect 10 122 766 128
<< labels >>
flabel comment s 176 403 176 403 0 FreeSans 300 0 0 0 S
flabel comment s 176 403 176 403 0 FreeSans 300 0 0 0 S
flabel comment s 282 403 282 403 0 FreeSans 300 0 0 0 S
flabel comment s 282 403 282 403 0 FreeSans 300 0 0 0 D
flabel comment s 388 403 388 403 0 FreeSans 300 0 0 0 S
flabel comment s 388 403 388 403 0 FreeSans 300 0 0 0 S
flabel comment s 494 403 494 403 0 FreeSans 300 0 0 0 S
flabel comment s 494 403 494 403 0 FreeSans 300 0 0 0 D
flabel comment s 600 403 600 403 0 FreeSans 300 0 0 0 S
flabel metal1 s 694 401 728 412 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal1 s 359 759 417 784 0 FreeSans 100 0 0 0 GATE
port 2 nsew
flabel metal1 s 359 17 417 42 0 FreeSans 100 0 0 0 GATE
port 2 nsew
flabel metal1 s 48 399 82 410 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal2 s 50 520 65 586 0 FreeSans 100 0 0 0 DRAIN
port 3 nsew
flabel metal2 s 59 205 73 268 0 FreeSans 100 0 0 0 SOURCE
port 4 nsew
<< properties >>
string GDS_END 9508088
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 9492266
<< end >>
