magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 2466 897
<< pwell >>
rect 2134 289 2396 317
rect 4 223 426 237
rect 1153 223 1435 289
rect 1862 223 2396 289
rect 4 43 2396 223
rect -26 -43 2426 43
<< locali >>
rect 108 381 174 515
rect 319 311 494 350
rect 2312 437 2378 747
rect 2328 137 2378 437
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2400 831
rect 108 735 298 741
rect 22 345 72 713
rect 108 701 114 735
rect 148 701 186 735
rect 220 701 258 735
rect 292 701 298 735
rect 444 735 494 741
rect 108 551 298 701
rect 334 523 400 713
rect 444 701 450 735
rect 484 701 494 735
rect 444 559 494 701
rect 1014 737 1204 747
rect 1014 703 1020 737
rect 1054 703 1092 737
rect 1126 703 1164 737
rect 1198 703 1204 737
rect 1014 697 1204 703
rect 530 661 736 695
rect 530 523 564 661
rect 702 627 1531 661
rect 334 489 564 523
rect 600 456 666 625
rect 702 492 768 627
rect 811 535 877 591
rect 1294 551 1461 591
rect 233 386 564 445
rect 600 422 807 456
rect 233 345 283 386
rect 530 352 737 386
rect 22 311 283 345
rect 22 119 76 311
rect 338 241 623 275
rect 686 241 737 352
rect 112 113 302 219
rect 338 119 404 241
rect 112 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 302 113
rect 112 73 302 79
rect 440 113 553 205
rect 440 79 443 113
rect 477 79 515 113
rect 549 79 553 113
rect 440 73 553 79
rect 589 87 623 241
rect 773 205 807 422
rect 659 123 807 205
rect 843 339 877 535
rect 913 477 1391 511
rect 913 377 978 477
rect 1341 445 1391 477
rect 1087 409 1153 441
rect 1427 409 1461 551
rect 1087 375 1461 409
rect 1497 503 1531 627
rect 1567 573 1617 747
rect 1763 735 1953 747
rect 1763 701 1769 735
rect 1803 701 1841 735
rect 1875 701 1913 735
rect 1947 701 1953 735
rect 1567 539 1720 573
rect 1763 539 1953 701
rect 1497 445 1650 503
rect 1686 489 1720 539
rect 1686 455 2007 489
rect 843 305 1269 339
rect 843 123 909 305
rect 945 235 1311 269
rect 945 87 1011 235
rect 589 53 1011 87
rect 1051 113 1241 199
rect 1051 79 1057 113
rect 1091 79 1129 113
rect 1163 79 1201 113
rect 1235 79 1241 113
rect 1051 73 1241 79
rect 1277 87 1311 235
rect 1347 123 1413 375
rect 1497 289 1531 445
rect 1456 225 1531 289
rect 1456 87 1490 225
rect 1686 205 1720 455
rect 1800 319 1866 403
rect 1941 355 2007 455
rect 2043 401 2109 747
rect 2145 735 2263 747
rect 2145 701 2151 735
rect 2185 701 2223 735
rect 2257 701 2263 735
rect 2145 439 2263 701
rect 2043 335 2292 401
rect 2043 319 2102 335
rect 1800 285 2102 319
rect 1567 189 1720 205
rect 1526 171 1720 189
rect 1526 105 1601 171
rect 1756 113 1946 249
rect 1277 53 1490 87
rect 1756 79 1762 113
rect 1796 79 1834 113
rect 1868 79 1906 113
rect 1940 79 1946 113
rect 2036 105 2102 285
rect 2138 113 2256 299
rect 1756 73 1946 79
rect 2138 79 2144 113
rect 2178 79 2216 113
rect 2250 79 2256 113
rect 2138 73 2256 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 114 701 148 735
rect 186 701 220 735
rect 258 701 292 735
rect 450 701 484 735
rect 1020 703 1054 737
rect 1092 703 1126 737
rect 1164 703 1198 737
rect 118 79 152 113
rect 190 79 224 113
rect 262 79 296 113
rect 443 79 477 113
rect 515 79 549 113
rect 1769 701 1803 735
rect 1841 701 1875 735
rect 1913 701 1947 735
rect 1057 79 1091 113
rect 1129 79 1163 113
rect 1201 79 1235 113
rect 2151 701 2185 735
rect 2223 701 2257 735
rect 1762 79 1796 113
rect 1834 79 1868 113
rect 1906 79 1940 113
rect 2144 79 2178 113
rect 2216 79 2250 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 831 2400 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2400 831
rect 0 791 2400 797
rect 0 737 2400 763
rect 0 735 1020 737
rect 0 701 114 735
rect 148 701 186 735
rect 220 701 258 735
rect 292 701 450 735
rect 484 703 1020 735
rect 1054 703 1092 737
rect 1126 703 1164 737
rect 1198 735 2400 737
rect 1198 703 1769 735
rect 484 701 1769 703
rect 1803 701 1841 735
rect 1875 701 1913 735
rect 1947 701 2151 735
rect 2185 701 2223 735
rect 2257 701 2400 735
rect 0 689 2400 701
rect 0 113 2400 125
rect 0 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 443 113
rect 477 79 515 113
rect 549 79 1057 113
rect 1091 79 1129 113
rect 1163 79 1201 113
rect 1235 79 1762 113
rect 1796 79 1834 113
rect 1868 79 1906 113
rect 1940 79 2144 113
rect 2178 79 2216 113
rect 2250 79 2400 113
rect 0 51 2400 79
rect 0 17 2400 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -23 2400 -17
<< labels >>
rlabel locali s 108 381 174 515 6 CLK
port 1 nsew clock input
rlabel locali s 319 311 494 350 6 D
port 2 nsew signal input
rlabel metal1 s 0 51 2400 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 2400 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 2426 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 43 2396 223 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1862 223 2396 289 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1153 223 1435 289 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 223 426 237 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 2134 289 2396 317 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 2400 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 2466 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 2400 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 2328 137 2378 437 6 Q
port 7 nsew signal output
rlabel locali s 2312 437 2378 747 6 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2400 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1154778
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 1130742
<< end >>
