magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 8 0 9 8 6 C0
port 1 nsew
rlabel  s 7 4 7 8 6 C0
port 1 nsew
rlabel  s 7 0 7 3 6 C0
port 1 nsew
rlabel  s 5 4 6 8 6 C0
port 1 nsew
rlabel  s 5 0 6 3 6 C0
port 1 nsew
rlabel  s 4 4 4 8 6 C0
port 1 nsew
rlabel  s 4 0 4 3 6 C0
port 1 nsew
rlabel  s 3 4 3 8 6 C0
port 1 nsew
rlabel  s 3 0 3 3 6 C0
port 1 nsew
rlabel  s 1 4 2 8 6 C0
port 1 nsew
rlabel  s 1 0 2 3 6 C0
port 1 nsew
rlabel  s 0 8 9 8 6 C0
port 1 nsew
rlabel  s 0 0 0 8 4 C0
port 1 nsew
rlabel  s 0 0 9 0 8 C0
port 1 nsew
rlabel  s 8 4 8 7 6 C1
port 2 nsew
rlabel  s 8 1 8 4 6 C1
port 2 nsew
rlabel  s 6 4 7 7 6 C1
port 2 nsew
rlabel  s 6 1 7 4 6 C1
port 2 nsew
rlabel  s 5 4 5 7 6 C1
port 2 nsew
rlabel  s 5 1 5 4 6 C1
port 2 nsew
rlabel  s 3 4 4 7 6 C1
port 2 nsew
rlabel  s 3 1 4 4 6 C1
port 2 nsew
rlabel  s 2 4 2 7 6 C1
port 2 nsew
rlabel  s 2 1 2 4 6 C1
port 2 nsew
rlabel  s 1 4 1 7 6 C1
port 2 nsew
rlabel  s 1 4 8 4 6 C1
port 2 nsew
rlabel  s 1 1 1 4 6 C1
port 2 nsew
rlabel r s 0 0 9 8 6 MET5
port 3 nsew
rlabel metal_blue s 4 4 5 4 6 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 9 8
string LEFview TRUE
<< end >>
