magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 8 2 8 8 6 B
port 1 nsew
rlabel  s 2 8 8 8 6 B
port 1 nsew
rlabel  s 2 6 2 8 6 B
port 1 nsew
rlabel  s 2 2 2 4 6 B
port 1 nsew
rlabel  s 2 2 8 2 6 B
port 1 nsew
rlabel  s 9 1 9 9 6 C
port 2 nsew
rlabel  s 1 9 9 9 6 C
port 2 nsew
rlabel  s 1 1 1 9 6 C
port 2 nsew
rlabel  s 1 1 9 1 6 C
port 2 nsew
rlabel  s 1 4 2 5 6 E
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 10 10
string LEFview TRUE
<< end >>
