magic
tech sky130B
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1663361622
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_1
timestamp 1663361622
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_2
timestamp 1663361622
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1663361622
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_1
timestamp 1663361622
transform 1 0 648 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 35265818
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 35263018
<< end >>
