magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 4 4 4 4 6 C0
port 1 nsew
rlabel  s 4 3 4 4 6 C0
port 1 nsew
rlabel  s 4 3 4 3 6 C0
port 1 nsew
rlabel  s 4 3 4 3 6 C0
port 1 nsew
rlabel  s 4 2 4 2 6 C0
port 1 nsew
rlabel  s 4 1 4 2 6 C0
port 1 nsew
rlabel  s 4 1 4 1 6 C0
port 1 nsew
rlabel  s 4 0 4 1 8 C0
port 1 nsew
rlabel  s 2 4 4 5 6 C0
port 1 nsew
rlabel  s 2 4 4 4 6 C0
port 1 nsew
rlabel  s 2 3 4 3 6 C0
port 1 nsew
rlabel  s 2 3 4 3 6 C0
port 1 nsew
rlabel  s 2 2 4 2 6 C0
port 1 nsew
rlabel  s 2 1 4 1 6 C0
port 1 nsew
rlabel  s 2 1 4 1 6 C0
port 1 nsew
rlabel  s 2 0 4 0 8 C0
port 1 nsew
rlabel  s 0 4 2 5 6 C0
port 1 nsew
rlabel  s 0 4 0 4 4 C0
port 1 nsew
rlabel  s 0 4 2 4 6 C0
port 1 nsew
rlabel  s 0 3 0 4 4 C0
port 1 nsew
rlabel  s 0 3 2 3 6 C0
port 1 nsew
rlabel  s 0 3 0 3 4 C0
port 1 nsew
rlabel  s 0 3 2 3 6 C0
port 1 nsew
rlabel  s 0 3 0 3 4 C0
port 1 nsew
rlabel  s 0 2 0 2 4 C0
port 1 nsew
rlabel  s 0 2 2 2 6 C0
port 1 nsew
rlabel  s 0 1 0 2 4 C0
port 1 nsew
rlabel  s 0 1 2 1 6 C0
port 1 nsew
rlabel  s 0 1 0 1 4 C0
port 1 nsew
rlabel  s 0 1 2 1 6 C0
port 1 nsew
rlabel  s 0 0 0 1 2 C0
port 1 nsew
rlabel  s 0 0 2 0 8 C0
port 1 nsew
rlabel  s 2 4 2 5 6 C1
port 2 nsew
rlabel  s 2 4 2 4 6 C1
port 2 nsew
rlabel  s 2 3 2 3 6 C1
port 2 nsew
rlabel  s 2 2 2 3 6 C1
port 2 nsew
rlabel  s 2 2 2 2 6 C1
port 2 nsew
rlabel  s 2 1 2 2 6 C1
port 2 nsew
rlabel  s 2 1 2 1 6 C1
port 2 nsew
rlabel  s 2 0 2 0 8 C1
port 2 nsew
rlabel  s 0 4 4 4 6 C1
port 2 nsew
rlabel  s 0 3 4 4 6 C1
port 2 nsew
rlabel  s 0 3 4 3 6 C1
port 2 nsew
rlabel  s 0 2 4 2 6 C1
port 2 nsew
rlabel  s 0 1 4 1 6 C1
port 2 nsew
rlabel  s 0 0 4 1 8 C1
port 2 nsew
rlabel  s 0 2 4 2 6 C1
port 2 nsew
rlabel  s 0 0 4 5 6 MET3
port 4 nsew
rlabel metal_blue s 2 2 2 2 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 4 5
string LEFview TRUE
<< end >>
