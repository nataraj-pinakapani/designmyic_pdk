magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 53 0 56 1 8 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 57 1 60 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 48 0 51 1 8 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 52 1 55 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 9 0 13 1 8 VCCD
port 3 nsew signal bidirectional
rlabel  s 0 13 1 17 4 VCCD
port 3 nsew signal bidirectional
rlabel  s 9 0 14 1 8 VCCD
port 3 nsew signal bidirectional
rlabel  s 0 13 1 17 4 VCCD
port 3 nsew signal bidirectional
rlabel  s 2 0 7 1 8 VCCHIB
port 4 nsew signal bidirectional
rlabel  s 0 6 1 11 4 VCCHIB
port 4 nsew signal bidirectional
rlabel  s 2 0 7 1 8 VCCHIB
port 4 nsew signal bidirectional
rlabel  s 0 6 1 11 4 VCCHIB
port 4 nsew signal bidirectional
rlabel  s 15 0 18 1 8 VDDA
port 5 nsew signal bidirectional
rlabel  s 0 19 1 22 4 VDDA
port 5 nsew signal bidirectional
rlabel  s 15 0 18 1 8 VDDA
port 5 nsew signal bidirectional
rlabel  s 0 19 1 22 4 VDDA
port 5 nsew signal bidirectional
rlabel  s 70 0 95 1 8 VDDIO
port 6 nsew signal bidirectional
rlabel  s 20 0 24 1 8 VDDIO
port 6 nsew signal bidirectional
rlabel  s 0 74 1 99 4 VDDIO
port 6 nsew signal bidirectional
rlabel  s 0 24 1 28 4 VDDIO
port 6 nsew signal bidirectional
rlabel  s 70 0 95 1 8 VDDIO
port 6 nsew signal bidirectional
rlabel  s 20 0 24 1 8 VDDIO
port 6 nsew signal bidirectional
rlabel  s 0 74 1 99 4 VDDIO
port 6 nsew signal bidirectional
rlabel  s 0 23 1 28 4 VDDIO
port 6 nsew signal bidirectional
rlabel  s 64 0 68 1 8 VDDIO_Q
port 7 nsew signal bidirectional
rlabel  s 0 68 1 72 4 VDDIO_Q
port 7 nsew signal bidirectional
rlabel  s 64 0 69 1 8 VDDIO_Q
port 7 nsew signal bidirectional
rlabel  s 0 68 1 72 4 VDDIO_Q
port 7 nsew signal bidirectional
rlabel  s 48 0 57 1 8 VSSA
port 8 nsew signal bidirectional
rlabel  s 37 0 40 1 8 VSSA
port 8 nsew signal bidirectional
rlabel  s 0 51 1 60 4 VSSA
port 8 nsew signal bidirectional
rlabel  s 0 41 1 44 4 VSSA
port 8 nsew signal bidirectional
rlabel  s 56 0 57 1 8 VSSA
port 8 nsew signal bidirectional
rlabel  s 52 0 53 1 8 VSSA
port 8 nsew signal bidirectional
rlabel  s 48 0 48 1 8 VSSA
port 8 nsew signal bidirectional
rlabel  s 37 0 40 1 8 VSSA
port 8 nsew signal bidirectional
rlabel  s 0 60 1 60 4 VSSA
port 8 nsew signal bidirectional
rlabel  s 0 55 1 56 4 VSSA
port 8 nsew signal bidirectional
rlabel  s 0 51 1 52 4 VSSA
port 8 nsew signal bidirectional
rlabel  s 0 40 1 44 4 VSSA
port 8 nsew signal bidirectional
rlabel  s 42 0 46 1 8 VSSD
port 9 nsew signal bidirectional
rlabel  s 0 45 1 50 4 VSSD
port 9 nsew signal bidirectional
rlabel  s 42 0 46 1 8 VSSD
port 9 nsew signal bidirectional
rlabel  s 0 45 1 50 4 VSSD
port 9 nsew signal bidirectional
rlabel  s 0 179 1 204 4 VSSIO
port 10 nsew signal bidirectional
rlabel  s 0 30 1 34 4 VSSIO
port 10 nsew signal bidirectional
rlabel  s 176 0 200 1 8 VSSIO
port 10 nsew signal bidirectional
rlabel  s 26 0 30 1 8 VSSIO
port 10 nsew signal bidirectional
rlabel  s 0 30 1 34 4 VSSIO
port 10 nsew signal bidirectional
rlabel  s 0 179 1 204 4 VSSIO
port 10 nsew signal bidirectional
rlabel  s 176 0 200 1 8 VSSIO
port 10 nsew signal bidirectional
rlabel  s 26 0 30 1 8 VSSIO
port 10 nsew signal bidirectional
rlabel  s 58 0 63 1 8 VSSIO_Q
port 11 nsew signal bidirectional
rlabel  s 0 62 1 66 4 VSSIO_Q
port 11 nsew signal bidirectional
rlabel  s 58 0 63 1 8 VSSIO_Q
port 11 nsew signal bidirectional
rlabel  s 0 62 1 66 4 VSSIO_Q
port 11 nsew signal bidirectional
rlabel  s 32 0 35 1 8 VSWITCH
port 12 nsew signal bidirectional
rlabel  s 0 36 1 39 4 VSWITCH
port 12 nsew signal bidirectional
rlabel  s 32 0 35 1 8 VSWITCH
port 12 nsew signal bidirectional
rlabel  s 0 36 1 39 4 VSWITCH
port 12 nsew signal bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 200 204
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
