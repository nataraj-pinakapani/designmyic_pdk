magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 710 157 892 201
rect 1200 157 1741 203
rect 1 21 1741 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 446 47 476 119
rect 542 47 572 119
rect 640 47 670 131
rect 786 47 816 175
rect 887 47 917 119
rect 990 47 1020 119
rect 1085 47 1115 131
rect 1278 47 1308 177
rect 1373 47 1403 177
rect 1457 47 1487 177
rect 1544 47 1574 177
rect 1628 47 1658 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 413 381 497
rect 445 413 475 497
rect 538 413 568 497
rect 634 413 664 497
rect 766 347 796 497
rect 861 413 891 497
rect 945 413 975 497
rect 1062 413 1092 497
rect 1278 297 1308 497
rect 1373 297 1403 497
rect 1457 297 1487 497
rect 1544 297 1574 497
rect 1628 297 1658 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 131
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 131
rect 736 131 786 175
rect 590 119 640 131
rect 381 107 446 119
rect 381 73 394 107
rect 428 73 446 107
rect 381 47 446 73
rect 476 107 542 119
rect 476 73 496 107
rect 530 73 542 107
rect 476 47 542 73
rect 572 47 640 119
rect 670 101 786 131
rect 670 67 714 101
rect 748 67 786 101
rect 670 47 786 67
rect 816 119 866 175
rect 1226 164 1278 177
rect 1035 119 1085 131
rect 816 107 887 119
rect 816 73 832 107
rect 866 73 887 107
rect 816 47 887 73
rect 917 107 990 119
rect 917 73 944 107
rect 978 73 990 107
rect 917 47 990 73
rect 1020 47 1085 119
rect 1115 107 1172 131
rect 1115 73 1125 107
rect 1159 73 1172 107
rect 1115 47 1172 73
rect 1226 130 1234 164
rect 1268 130 1278 164
rect 1226 96 1278 130
rect 1226 62 1234 96
rect 1268 62 1278 96
rect 1226 47 1278 62
rect 1308 97 1373 177
rect 1308 63 1325 97
rect 1359 63 1373 97
rect 1308 47 1373 63
rect 1403 164 1457 177
rect 1403 130 1413 164
rect 1447 130 1457 164
rect 1403 96 1457 130
rect 1403 62 1413 96
rect 1447 62 1457 96
rect 1403 47 1457 62
rect 1487 96 1544 177
rect 1487 62 1499 96
rect 1533 62 1544 96
rect 1487 47 1544 62
rect 1574 164 1628 177
rect 1574 130 1584 164
rect 1618 130 1628 164
rect 1574 96 1628 130
rect 1574 62 1584 96
rect 1618 62 1628 96
rect 1574 47 1628 62
rect 1658 96 1715 177
rect 1658 62 1669 96
rect 1703 62 1715 96
rect 1658 47 1715 62
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 413 351 451
rect 381 472 445 497
rect 381 438 391 472
rect 425 438 445 472
rect 381 413 445 438
rect 475 472 538 497
rect 475 438 490 472
rect 524 438 538 472
rect 475 413 538 438
rect 568 413 634 497
rect 664 485 766 497
rect 664 451 722 485
rect 756 451 766 485
rect 664 417 766 451
rect 664 413 722 417
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 679 383 722 413
rect 756 383 766 417
rect 679 347 766 383
rect 796 477 861 497
rect 796 443 806 477
rect 840 443 861 477
rect 796 413 861 443
rect 891 467 945 497
rect 891 433 901 467
rect 935 433 945 467
rect 891 413 945 433
rect 975 413 1062 497
rect 1092 477 1150 497
rect 1092 443 1102 477
rect 1136 443 1150 477
rect 1092 413 1150 443
rect 1222 475 1278 497
rect 1222 441 1234 475
rect 1268 441 1278 475
rect 796 347 846 413
rect 1222 407 1278 441
rect 1222 373 1234 407
rect 1268 373 1278 407
rect 1222 339 1278 373
rect 1222 305 1234 339
rect 1268 305 1278 339
rect 1222 297 1278 305
rect 1308 489 1373 497
rect 1308 455 1325 489
rect 1359 455 1373 489
rect 1308 421 1373 455
rect 1308 387 1325 421
rect 1359 387 1373 421
rect 1308 297 1373 387
rect 1403 479 1457 497
rect 1403 445 1413 479
rect 1447 445 1457 479
rect 1403 411 1457 445
rect 1403 377 1413 411
rect 1447 377 1457 411
rect 1403 343 1457 377
rect 1403 309 1413 343
rect 1447 309 1457 343
rect 1403 297 1457 309
rect 1487 479 1544 497
rect 1487 445 1500 479
rect 1534 445 1544 479
rect 1487 411 1544 445
rect 1487 377 1500 411
rect 1534 377 1544 411
rect 1487 297 1544 377
rect 1574 479 1628 497
rect 1574 445 1584 479
rect 1618 445 1628 479
rect 1574 411 1628 445
rect 1574 377 1584 411
rect 1618 377 1628 411
rect 1574 343 1628 377
rect 1574 309 1584 343
rect 1618 309 1628 343
rect 1574 297 1628 309
rect 1658 479 1714 497
rect 1658 445 1668 479
rect 1702 445 1714 479
rect 1658 411 1714 445
rect 1658 377 1668 411
rect 1702 377 1714 411
rect 1658 297 1714 377
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 394 73 428 107
rect 496 73 530 107
rect 714 67 748 101
rect 832 73 866 107
rect 944 73 978 107
rect 1125 73 1159 107
rect 1234 130 1268 164
rect 1234 62 1268 96
rect 1325 63 1359 97
rect 1413 130 1447 164
rect 1413 62 1447 96
rect 1499 62 1533 96
rect 1584 130 1618 164
rect 1584 62 1618 96
rect 1669 62 1703 96
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 307 451 341 485
rect 391 438 425 472
rect 490 438 524 472
rect 722 451 756 485
rect 203 375 237 409
rect 722 383 756 417
rect 806 443 840 477
rect 901 433 935 467
rect 1102 443 1136 477
rect 1234 441 1268 475
rect 1234 373 1268 407
rect 1234 305 1268 339
rect 1325 455 1359 489
rect 1325 387 1359 421
rect 1413 445 1447 479
rect 1413 377 1447 411
rect 1413 309 1447 343
rect 1500 445 1534 479
rect 1500 377 1534 411
rect 1584 445 1618 479
rect 1584 377 1618 411
rect 1584 309 1618 343
rect 1668 445 1702 479
rect 1668 377 1702 411
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 445 497 475 523
rect 538 497 568 523
rect 634 497 664 523
rect 766 497 796 523
rect 861 497 891 523
rect 945 497 975 523
rect 1062 497 1092 523
rect 1278 497 1308 523
rect 1373 497 1403 523
rect 1457 497 1487 523
rect 1544 497 1574 523
rect 1628 497 1658 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 265 76 318
rect 163 274 193 363
rect 351 333 381 413
rect 445 375 475 413
rect 538 381 568 413
rect 22 249 76 265
rect 22 215 32 249
rect 66 215 76 249
rect 118 264 193 274
rect 300 317 381 333
rect 430 365 496 375
rect 430 331 446 365
rect 480 331 496 365
rect 430 321 496 331
rect 538 365 592 381
rect 538 331 548 365
rect 582 331 592 365
rect 300 283 310 317
rect 344 283 381 317
rect 300 267 381 283
rect 538 315 592 331
rect 538 279 568 315
rect 118 230 134 264
rect 168 230 193 264
rect 118 220 193 230
rect 22 199 76 215
rect 46 176 76 199
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 351 131 381 267
rect 446 249 568 279
rect 446 119 476 249
rect 634 213 664 413
rect 766 309 796 347
rect 861 315 891 413
rect 945 375 975 413
rect 944 365 1010 375
rect 944 331 960 365
rect 994 331 1010 365
rect 944 321 1010 331
rect 1062 366 1092 413
rect 1062 350 1140 366
rect 1062 316 1096 350
rect 1130 316 1140 350
rect 706 299 796 309
rect 706 265 722 299
rect 756 265 796 299
rect 706 255 796 265
rect 766 220 796 255
rect 848 299 902 315
rect 1062 300 1140 316
rect 848 265 858 299
rect 892 279 902 299
rect 892 265 1020 279
rect 848 249 1020 265
rect 518 191 572 207
rect 518 157 528 191
rect 562 157 572 191
rect 634 203 714 213
rect 634 183 664 203
rect 518 141 572 157
rect 542 119 572 141
rect 640 169 664 183
rect 698 169 714 203
rect 766 190 816 220
rect 786 175 816 190
rect 887 191 948 207
rect 640 159 714 169
rect 640 131 670 159
rect 887 157 904 191
rect 938 157 948 191
rect 887 141 948 157
rect 887 119 917 141
rect 990 119 1020 249
rect 1085 131 1115 300
rect 1278 265 1308 297
rect 1186 249 1308 265
rect 1186 215 1196 249
rect 1230 215 1308 249
rect 1186 199 1308 215
rect 1278 177 1308 199
rect 1373 265 1403 297
rect 1457 265 1487 297
rect 1544 265 1574 297
rect 1628 265 1658 297
rect 1373 249 1658 265
rect 1373 215 1394 249
rect 1428 215 1462 249
rect 1496 215 1530 249
rect 1564 215 1598 249
rect 1632 215 1658 249
rect 1373 199 1658 215
rect 1373 177 1403 199
rect 1457 177 1487 199
rect 1544 177 1574 199
rect 1628 177 1658 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 446 21 476 47
rect 542 21 572 47
rect 640 21 670 47
rect 786 21 816 47
rect 887 21 917 47
rect 990 21 1020 47
rect 1085 21 1115 47
rect 1278 21 1308 47
rect 1373 21 1403 47
rect 1457 21 1487 47
rect 1544 21 1574 47
rect 1628 21 1658 47
<< polycont >>
rect 32 215 66 249
rect 446 331 480 365
rect 548 331 582 365
rect 310 283 344 317
rect 134 230 168 264
rect 960 331 994 365
rect 1096 316 1130 350
rect 722 265 756 299
rect 858 265 892 299
rect 528 157 562 191
rect 664 169 698 203
rect 904 157 938 191
rect 1196 215 1230 249
rect 1394 215 1428 249
rect 1462 215 1496 249
rect 1530 215 1564 249
rect 1598 215 1632 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 203 409 248 443
rect 288 485 341 527
rect 288 451 307 485
rect 288 435 341 451
rect 378 472 425 488
rect 722 485 756 527
rect 378 438 391 472
rect 474 438 490 472
rect 524 438 688 472
rect 69 391 168 393
rect 69 375 122 391
rect 35 359 122 375
rect 156 357 168 391
rect 18 249 88 325
rect 18 215 32 249
rect 66 215 88 249
rect 18 195 88 215
rect 122 264 168 357
rect 122 230 134 264
rect 122 161 168 230
rect 35 127 168 161
rect 237 375 248 409
rect 203 187 248 375
rect 378 413 425 438
rect 288 317 344 333
rect 288 283 310 317
rect 288 213 344 283
rect 203 153 214 187
rect 35 119 69 127
rect 203 119 248 153
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 248 119
rect 203 69 248 85
rect 291 93 341 109
rect 103 17 169 59
rect 291 59 307 93
rect 378 107 412 413
rect 532 391 620 402
rect 446 365 494 381
rect 480 331 494 365
rect 532 365 586 391
rect 532 331 548 365
rect 582 357 586 365
rect 582 331 620 357
rect 446 207 494 331
rect 654 315 688 438
rect 722 417 756 451
rect 722 367 756 383
rect 790 477 840 493
rect 790 443 806 477
rect 1098 477 1141 527
rect 790 427 840 443
rect 885 433 901 467
rect 935 433 1062 467
rect 654 299 756 315
rect 654 297 722 299
rect 596 265 722 297
rect 596 263 756 265
rect 446 191 562 207
rect 446 187 528 191
rect 446 153 494 187
rect 528 153 562 157
rect 446 141 562 153
rect 596 107 630 263
rect 722 249 756 263
rect 664 213 698 219
rect 790 213 824 427
rect 858 391 896 393
rect 858 357 862 391
rect 858 299 896 357
rect 892 265 896 299
rect 858 249 896 265
rect 930 365 994 381
rect 930 331 960 365
rect 930 315 994 331
rect 664 203 824 213
rect 930 207 968 315
rect 698 169 824 203
rect 664 153 824 169
rect 378 73 394 107
rect 428 73 444 107
rect 480 73 496 107
rect 530 73 630 107
rect 680 101 754 117
rect 291 17 341 59
rect 680 67 714 101
rect 748 67 754 101
rect 790 107 824 153
rect 858 191 968 207
rect 858 187 904 191
rect 858 153 862 187
rect 896 157 904 187
rect 938 157 968 191
rect 896 153 968 157
rect 858 141 968 153
rect 1028 249 1062 433
rect 1098 443 1102 477
rect 1136 443 1141 477
rect 1098 427 1141 443
rect 1234 475 1268 491
rect 1234 407 1268 441
rect 1234 366 1268 373
rect 1325 489 1361 527
rect 1359 455 1361 489
rect 1500 479 1534 527
rect 1668 479 1702 527
rect 1325 421 1361 455
rect 1359 387 1361 421
rect 1325 371 1361 387
rect 1397 445 1413 479
rect 1447 445 1464 479
rect 1397 411 1464 445
rect 1397 377 1413 411
rect 1447 377 1464 411
rect 1096 350 1268 366
rect 1130 339 1268 350
rect 1130 316 1234 339
rect 1096 305 1234 316
rect 1397 343 1464 377
rect 1500 411 1534 445
rect 1500 361 1534 377
rect 1568 445 1584 479
rect 1618 445 1634 479
rect 1568 411 1634 445
rect 1568 377 1584 411
rect 1618 377 1634 411
rect 1268 305 1318 334
rect 1096 300 1318 305
rect 1284 249 1318 300
rect 1397 309 1413 343
rect 1447 327 1464 343
rect 1568 343 1634 377
rect 1668 411 1702 445
rect 1668 361 1702 377
rect 1568 327 1584 343
rect 1447 309 1584 327
rect 1618 327 1634 343
rect 1618 309 1731 327
rect 1397 293 1731 309
rect 1028 215 1196 249
rect 1230 215 1246 249
rect 1284 215 1394 249
rect 1428 215 1462 249
rect 1496 215 1530 249
rect 1564 215 1598 249
rect 1632 215 1648 249
rect 1028 107 1062 215
rect 1284 181 1318 215
rect 1218 164 1318 181
rect 1682 180 1731 293
rect 1218 130 1234 164
rect 1268 147 1318 164
rect 1397 164 1731 180
rect 1268 130 1290 147
rect 790 73 832 107
rect 866 73 882 107
rect 928 73 944 107
rect 978 73 1062 107
rect 1125 107 1159 123
rect 680 17 754 67
rect 1125 17 1159 73
rect 1218 96 1290 130
rect 1397 130 1413 164
rect 1447 146 1584 164
rect 1447 130 1464 146
rect 1218 62 1234 96
rect 1268 62 1290 96
rect 1218 59 1290 62
rect 1325 97 1359 113
rect 1325 17 1359 63
rect 1397 96 1464 130
rect 1568 130 1584 146
rect 1618 146 1731 164
rect 1618 130 1635 146
rect 1397 62 1413 96
rect 1447 62 1464 96
rect 1397 61 1464 62
rect 1499 96 1533 112
rect 1499 17 1533 62
rect 1568 96 1635 130
rect 1568 62 1584 96
rect 1618 62 1635 96
rect 1568 61 1635 62
rect 1669 96 1703 112
rect 1669 17 1703 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 122 357 156 391
rect 214 153 248 187
rect 586 357 620 391
rect 494 153 528 187
rect 862 357 896 391
rect 862 153 896 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 110 391 168 397
rect 110 357 122 391
rect 156 388 168 391
rect 574 391 632 397
rect 574 388 586 391
rect 156 360 586 388
rect 156 357 168 360
rect 110 351 168 357
rect 574 357 586 360
rect 620 388 632 391
rect 850 391 908 397
rect 850 388 862 391
rect 620 360 862 388
rect 620 357 632 360
rect 574 351 632 357
rect 850 357 862 360
rect 896 357 908 391
rect 850 351 908 357
rect 202 187 260 193
rect 202 153 214 187
rect 248 184 260 187
rect 482 187 540 193
rect 482 184 494 187
rect 248 156 494 184
rect 248 153 260 156
rect 202 147 260 153
rect 482 153 494 156
rect 528 184 540 187
rect 850 187 908 193
rect 850 184 862 187
rect 528 156 862 184
rect 528 153 540 156
rect 482 147 540 153
rect 850 153 862 156
rect 896 153 908 187
rect 850 147 908 153
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1409 85 1443 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1409 357 1443 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1409 425 1443 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 305 289 339 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 4 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 5 nsew
rlabel comment s 0 0 0 0 4 dfxtp_4
rlabel metal1 s 0 -48 1748 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_END 2723432
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 2709332
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 43.700 0.000 
<< end >>
