/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/lef/sky130_fd_sc_hvl/sky130_fd_sc_hvl.lef