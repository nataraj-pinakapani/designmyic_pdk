magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 1 1 2 1 6 C0
port 1 nsew
rlabel  s 1 0 2 1 8 C0
port 1 nsew
rlabel  s 1 1 2 2 6 C0
port 1 nsew
rlabel  s 1 0 2 0 8 C0
port 1 nsew
rlabel  s 0 1 1 2 4 C0
port 1 nsew
rlabel  s 0 1 0 1 4 C0
port 1 nsew
rlabel  s 0 0 0 1 2 C0
port 1 nsew
rlabel  s 0 0 1 0 2 C0
port 1 nsew
rlabel  s 1 1 1 2 6 C1
port 2 nsew
rlabel  s 1 1 1 1 6 C1
port 2 nsew
rlabel  s 1 1 1 1 6 C1
port 2 nsew
rlabel  s 1 0 1 0 8 C1
port 2 nsew
rlabel  s 0 1 1 1 4 C1
port 2 nsew
rlabel  s 0 0 1 1 2 C1
port 2 nsew
rlabel  s 0 1 2 1 6 C1
port 2 nsew
rlabel  s -1 -1 3 3 6 MET3
port 4 nsew
rlabel metal_blue s 1 1 1 1 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -1 -1 3 3
string LEFview TRUE
<< end >>
