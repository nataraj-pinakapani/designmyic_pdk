magic
tech sky130A
timestamp 1663361622
<< properties >>
string GDS_END 32427708
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 32427068
<< end >>
