magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 3 2 3 3 6 DRAIN
port 1 nsew
rlabel  s 2 2 3 3 6 DRAIN
port 1 nsew
rlabel  s 1 2 2 3 6 DRAIN
port 1 nsew
rlabel  s 1 3 3 3 6 DRAIN
port 1 nsew
rlabel  s 1 2 1 3 6 DRAIN
port 1 nsew
rlabel  s 1 3 3 4 6 GATE
port 2 nsew
rlabel  s 4 0 4 3 6 SOURCE
port 3 nsew
rlabel  s 3 0 3 3 6 SOURCE
port 3 nsew
rlabel  s 2 0 2 3 6 SOURCE
port 3 nsew
rlabel  s 1 0 1 3 6 SOURCE
port 3 nsew
rlabel  s 0 0 0 3 4 SOURCE
port 3 nsew
rlabel  s 0 0 4 0 8 SOURCE
port 3 nsew
rlabel metal_blue s 0 3 0 3 4 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 4 4
string LEFview TRUE
<< end >>
