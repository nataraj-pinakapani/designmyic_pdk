/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/fixed_devices/sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p15_fail.cdl