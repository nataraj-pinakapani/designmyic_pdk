magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 4 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 4 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 9 nsew power bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 9 nsew power bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string LEFclass PAD SPACER
string FIXED_BBOX 0 0 1 198
string LEFview TRUE
<< end >>
