magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 835 157 1471 203
rect 1 21 1471 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 352 47 382 131
rect 436 47 466 131
rect 544 47 574 119
rect 630 47 660 119
rect 725 47 755 131
rect 913 47 943 177
rect 997 47 1027 177
rect 1093 47 1123 177
rect 1184 47 1214 177
rect 1271 47 1301 177
rect 1363 47 1393 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 352 369 382 497
rect 436 369 466 497
rect 532 413 562 497
rect 653 413 683 497
rect 725 413 755 497
rect 913 297 943 497
rect 997 297 1027 497
rect 1093 297 1123 497
rect 1184 297 1214 497
rect 1271 297 1301 497
rect 1363 297 1393 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 300 119 352 131
rect 300 85 308 119
rect 342 85 352 119
rect 300 47 352 85
rect 382 89 436 131
rect 382 55 392 89
rect 426 55 436 89
rect 382 47 436 55
rect 466 119 516 131
rect 861 165 913 177
rect 861 131 869 165
rect 903 131 913 165
rect 675 119 725 131
rect 466 47 544 119
rect 574 107 630 119
rect 574 73 585 107
rect 619 73 630 107
rect 574 47 630 73
rect 660 47 725 119
rect 755 106 807 131
rect 755 72 765 106
rect 799 72 807 106
rect 755 47 807 72
rect 861 97 913 131
rect 861 63 869 97
rect 903 63 913 97
rect 861 47 913 63
rect 943 47 997 177
rect 1027 89 1093 177
rect 1027 55 1038 89
rect 1072 55 1093 89
rect 1027 47 1093 55
rect 1123 89 1184 177
rect 1123 55 1138 89
rect 1172 55 1184 89
rect 1123 47 1184 55
rect 1214 93 1271 177
rect 1214 59 1227 93
rect 1261 59 1271 93
rect 1214 47 1271 59
rect 1301 115 1363 177
rect 1301 81 1315 115
rect 1349 81 1363 115
rect 1301 47 1363 81
rect 1393 93 1445 177
rect 1393 59 1403 93
rect 1437 59 1445 93
rect 1393 47 1445 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 300 483 352 497
rect 300 449 308 483
rect 342 449 352 483
rect 300 415 352 449
rect 300 381 308 415
rect 342 381 352 415
rect 300 369 352 381
rect 382 485 436 497
rect 382 451 392 485
rect 426 451 436 485
rect 382 417 436 451
rect 382 383 392 417
rect 426 383 436 417
rect 382 369 436 383
rect 466 413 532 497
rect 562 485 653 497
rect 562 451 597 485
rect 631 451 653 485
rect 562 413 653 451
rect 683 413 725 497
rect 755 477 807 497
rect 755 443 765 477
rect 799 443 807 477
rect 755 413 807 443
rect 861 485 913 497
rect 861 451 869 485
rect 903 451 913 485
rect 466 369 516 413
rect 861 297 913 451
rect 943 471 997 497
rect 943 437 953 471
rect 987 437 997 471
rect 943 368 997 437
rect 943 334 953 368
rect 987 334 997 368
rect 943 297 997 334
rect 1027 489 1093 497
rect 1027 455 1043 489
rect 1077 455 1093 489
rect 1027 421 1093 455
rect 1027 387 1043 421
rect 1077 387 1093 421
rect 1027 297 1093 387
rect 1123 477 1184 497
rect 1123 443 1136 477
rect 1170 443 1184 477
rect 1123 297 1184 443
rect 1214 485 1271 497
rect 1214 451 1227 485
rect 1261 451 1271 485
rect 1214 417 1271 451
rect 1214 383 1227 417
rect 1261 383 1271 417
rect 1214 349 1271 383
rect 1214 315 1227 349
rect 1261 315 1271 349
rect 1214 297 1271 315
rect 1301 477 1363 497
rect 1301 443 1315 477
rect 1349 443 1363 477
rect 1301 409 1363 443
rect 1301 375 1315 409
rect 1349 375 1363 409
rect 1301 297 1363 375
rect 1393 485 1445 497
rect 1393 451 1403 485
rect 1437 451 1445 485
rect 1393 417 1445 451
rect 1393 383 1403 417
rect 1437 383 1445 417
rect 1393 349 1445 383
rect 1393 315 1403 349
rect 1437 315 1445 349
rect 1393 297 1445 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 308 85 342 119
rect 392 55 426 89
rect 869 131 903 165
rect 585 73 619 107
rect 765 72 799 106
rect 869 63 903 97
rect 1038 55 1072 89
rect 1138 55 1172 89
rect 1227 59 1261 93
rect 1315 81 1349 115
rect 1403 59 1437 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 308 449 342 483
rect 308 381 342 415
rect 392 451 426 485
rect 392 383 426 417
rect 597 451 631 485
rect 765 443 799 477
rect 869 451 903 485
rect 953 437 987 471
rect 953 334 987 368
rect 1043 455 1077 489
rect 1043 387 1077 421
rect 1136 443 1170 477
rect 1227 451 1261 485
rect 1227 383 1261 417
rect 1227 315 1261 349
rect 1315 443 1349 477
rect 1315 375 1349 409
rect 1403 451 1437 485
rect 1403 383 1437 417
rect 1403 315 1437 349
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 352 497 382 523
rect 436 497 466 523
rect 532 497 562 523
rect 653 497 683 523
rect 725 497 755 523
rect 913 497 943 523
rect 997 497 1027 523
rect 1093 497 1123 523
rect 1184 497 1214 523
rect 1271 497 1301 523
rect 1363 497 1393 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 352 241 382 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 299 225 382 241
rect 299 191 309 225
rect 343 191 382 225
rect 436 219 466 369
rect 532 337 562 413
rect 653 375 683 413
rect 508 321 562 337
rect 604 365 683 375
rect 604 331 620 365
rect 654 331 683 365
rect 604 321 683 331
rect 725 373 755 413
rect 725 357 813 373
rect 725 323 769 357
rect 803 323 813 357
rect 508 287 518 321
rect 552 287 562 321
rect 508 279 562 287
rect 725 307 813 323
rect 508 271 660 279
rect 532 249 660 271
rect 299 175 382 191
rect 352 131 382 175
rect 425 203 479 219
rect 425 169 435 203
rect 469 169 479 203
rect 425 153 479 169
rect 534 191 588 207
rect 534 157 544 191
rect 578 157 588 191
rect 436 131 466 153
rect 534 141 588 157
rect 544 119 574 141
rect 630 119 660 249
rect 725 131 755 307
rect 913 259 943 297
rect 997 265 1027 297
rect 1093 265 1123 297
rect 1184 265 1214 297
rect 1271 265 1301 297
rect 1363 265 1393 297
rect 797 249 943 259
rect 797 215 813 249
rect 847 215 943 249
rect 797 205 943 215
rect 913 177 943 205
rect 985 249 1039 265
rect 985 215 995 249
rect 1029 215 1039 249
rect 985 199 1039 215
rect 1081 249 1393 265
rect 1081 215 1091 249
rect 1125 215 1393 249
rect 1081 199 1393 215
rect 997 177 1027 199
rect 1093 177 1123 199
rect 1184 177 1214 199
rect 1271 177 1301 199
rect 1363 177 1393 199
rect 79 21 109 47
rect 163 21 193 47
rect 352 21 382 47
rect 436 21 466 47
rect 544 21 574 47
rect 630 21 660 47
rect 725 21 755 47
rect 913 21 943 47
rect 997 21 1027 47
rect 1093 21 1123 47
rect 1184 21 1214 47
rect 1271 21 1301 47
rect 1363 21 1393 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 309 191 343 225
rect 620 331 654 365
rect 769 323 803 357
rect 518 287 552 321
rect 435 169 469 203
rect 544 157 578 191
rect 813 215 847 249
rect 995 215 1029 249
rect 1091 215 1125 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 392 485 455 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 292 449 308 483
rect 342 449 358 483
rect 292 415 358 449
rect 292 381 308 415
rect 342 381 358 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 292 333 358 381
rect 426 451 455 485
rect 581 451 597 485
rect 631 451 731 485
rect 392 417 455 451
rect 426 383 455 417
rect 392 367 455 383
rect 586 391 654 399
rect 586 357 587 391
rect 621 365 654 391
rect 292 299 429 333
rect 293 225 359 265
rect 293 191 309 225
rect 343 191 359 225
rect 395 219 429 299
rect 495 323 552 337
rect 529 321 552 323
rect 495 287 518 289
rect 495 271 552 287
rect 586 331 620 357
rect 586 315 654 331
rect 395 203 469 219
rect 586 207 620 315
rect 697 265 731 451
rect 765 477 823 527
rect 799 443 823 477
rect 765 427 823 443
rect 861 485 917 527
rect 861 451 869 485
rect 903 451 917 485
rect 861 427 917 451
rect 951 471 989 493
rect 951 437 953 471
rect 987 437 989 471
rect 951 373 989 437
rect 1023 489 1097 527
rect 1023 455 1043 489
rect 1077 455 1097 489
rect 1023 421 1097 455
rect 1023 387 1043 421
rect 1077 387 1097 421
rect 1023 375 1097 387
rect 1136 477 1193 493
rect 1170 443 1193 477
rect 1136 375 1193 443
rect 765 368 989 373
rect 765 357 953 368
rect 765 323 769 357
rect 803 334 953 357
rect 987 341 989 368
rect 987 334 1125 341
rect 803 323 1125 334
rect 765 307 1125 323
rect 697 249 847 265
rect 697 233 813 249
rect 395 169 435 203
rect 395 157 469 169
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 308 153 469 157
rect 544 191 620 207
rect 578 157 620 191
rect 308 123 429 153
rect 544 141 620 157
rect 667 215 813 233
rect 667 199 847 215
rect 901 249 1029 265
rect 901 215 995 249
rect 901 199 1029 215
rect 1091 249 1125 307
rect 308 119 342 123
rect 667 107 701 199
rect 1091 165 1125 215
rect 308 69 342 85
rect 103 17 169 59
rect 376 55 392 89
rect 426 55 442 89
rect 569 73 585 107
rect 619 73 701 107
rect 853 131 869 165
rect 903 131 1125 165
rect 1159 265 1193 375
rect 1227 485 1281 527
rect 1261 451 1281 485
rect 1227 417 1281 451
rect 1261 383 1281 417
rect 1227 349 1281 383
rect 1261 315 1281 349
rect 1227 299 1281 315
rect 1315 477 1355 493
rect 1349 443 1355 477
rect 1315 409 1355 443
rect 1349 375 1355 409
rect 1315 265 1355 375
rect 1389 485 1455 527
rect 1389 451 1403 485
rect 1437 451 1455 485
rect 1389 417 1455 451
rect 1389 383 1403 417
rect 1437 383 1455 417
rect 1389 349 1455 383
rect 1389 315 1403 349
rect 1437 315 1455 349
rect 1389 299 1455 315
rect 1159 153 1455 265
rect 376 17 442 55
rect 749 72 765 106
rect 799 72 815 106
rect 749 17 815 72
rect 853 97 919 131
rect 1159 97 1193 153
rect 853 63 869 97
rect 903 63 919 97
rect 853 51 919 63
rect 1020 89 1088 97
rect 1020 55 1038 89
rect 1072 55 1088 89
rect 1020 17 1088 55
rect 1122 89 1193 97
rect 1122 55 1138 89
rect 1172 55 1193 89
rect 1122 51 1193 55
rect 1227 93 1281 119
rect 1261 59 1281 93
rect 1227 17 1281 59
rect 1315 115 1355 153
rect 1349 81 1355 115
rect 1315 51 1355 81
rect 1389 93 1455 119
rect 1389 59 1403 93
rect 1437 59 1455 93
rect 1389 17 1455 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 587 365 621 391
rect 587 357 620 365
rect 620 357 621 365
rect 495 321 529 323
rect 495 289 518 321
rect 518 289 529 321
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 575 391 633 397
rect 575 388 587 391
rect 248 360 587 388
rect 248 357 260 360
rect 202 351 260 357
rect 575 357 587 360
rect 621 357 633 391
rect 575 351 633 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 483 323 541 329
rect 483 320 495 323
rect 156 292 495 320
rect 156 289 168 292
rect 110 283 168 289
rect 483 289 495 292
rect 529 289 541 323
rect 483 283 541 289
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1235 153 1269 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1235 221 1269 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1419 153 1453 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1419 221 1453 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1327 221 1361 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 959 221 993 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1143 425 1177 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1327 153 1361 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 311 221 345 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 0 496 1472 592 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 dlrtp_4
rlabel metal1 s 0 -48 1472 48 1 VGND
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 2810794
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 2798072
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
