magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 6 21 827 203
rect 28 -17 62 21
<< scnmos >>
rect 84 47 114 177
rect 190 47 220 177
rect 274 47 304 177
rect 358 47 388 177
rect 464 47 494 177
rect 548 47 578 177
rect 632 47 662 177
rect 716 47 746 177
<< scpmoshvt >>
rect 84 297 114 497
rect 190 297 220 497
rect 274 297 304 497
rect 358 297 388 497
rect 464 297 494 497
rect 548 297 578 497
rect 632 297 662 497
rect 716 297 746 497
<< ndiff >>
rect 32 101 84 177
rect 32 67 40 101
rect 74 67 84 101
rect 32 47 84 67
rect 114 115 190 177
rect 114 81 140 115
rect 174 81 190 115
rect 114 47 190 81
rect 220 97 274 177
rect 220 63 230 97
rect 264 63 274 97
rect 220 47 274 63
rect 304 115 358 177
rect 304 81 314 115
rect 348 81 358 115
rect 304 47 358 81
rect 388 97 464 177
rect 388 63 418 97
rect 452 63 464 97
rect 388 47 464 63
rect 494 114 548 177
rect 494 80 504 114
rect 538 80 548 114
rect 494 47 548 80
rect 578 95 632 177
rect 578 61 588 95
rect 622 61 632 95
rect 578 47 632 61
rect 662 163 716 177
rect 662 129 672 163
rect 706 129 716 163
rect 662 95 716 129
rect 662 61 672 95
rect 706 61 716 95
rect 662 47 716 61
rect 746 95 801 177
rect 746 61 756 95
rect 790 61 801 95
rect 746 47 801 61
<< pdiff >>
rect 32 485 84 497
rect 32 451 40 485
rect 74 451 84 485
rect 32 417 84 451
rect 32 383 40 417
rect 74 383 84 417
rect 32 349 84 383
rect 32 315 40 349
rect 74 315 84 349
rect 32 297 84 315
rect 114 297 190 497
rect 220 297 274 497
rect 304 297 358 497
rect 388 477 464 497
rect 388 443 409 477
rect 443 443 464 477
rect 388 409 464 443
rect 388 375 409 409
rect 443 375 464 409
rect 388 297 464 375
rect 494 477 548 497
rect 494 443 504 477
rect 538 443 548 477
rect 494 409 548 443
rect 494 375 504 409
rect 538 375 548 409
rect 494 341 548 375
rect 494 307 504 341
rect 538 307 548 341
rect 494 297 548 307
rect 578 477 632 497
rect 578 443 588 477
rect 622 443 632 477
rect 578 409 632 443
rect 578 375 588 409
rect 622 375 632 409
rect 578 297 632 375
rect 662 477 716 497
rect 662 443 672 477
rect 706 443 716 477
rect 662 409 716 443
rect 662 375 672 409
rect 706 375 716 409
rect 662 341 716 375
rect 662 307 672 341
rect 706 307 716 341
rect 662 297 716 307
rect 746 477 800 497
rect 746 443 756 477
rect 790 443 800 477
rect 746 409 800 443
rect 746 375 756 409
rect 790 375 800 409
rect 746 297 800 375
<< ndiffc >>
rect 40 67 74 101
rect 140 81 174 115
rect 230 63 264 97
rect 314 81 348 115
rect 418 63 452 97
rect 504 80 538 114
rect 588 61 622 95
rect 672 129 706 163
rect 672 61 706 95
rect 756 61 790 95
<< pdiffc >>
rect 40 451 74 485
rect 40 383 74 417
rect 40 315 74 349
rect 409 443 443 477
rect 409 375 443 409
rect 504 443 538 477
rect 504 375 538 409
rect 504 307 538 341
rect 588 443 622 477
rect 588 375 622 409
rect 672 443 706 477
rect 672 375 706 409
rect 672 307 706 341
rect 756 443 790 477
rect 756 375 790 409
<< poly >>
rect 84 497 114 523
rect 190 497 220 523
rect 274 497 304 523
rect 358 497 388 523
rect 464 497 494 523
rect 548 497 578 523
rect 632 497 662 523
rect 716 497 746 523
rect 84 265 114 297
rect 190 265 220 297
rect 274 265 304 297
rect 358 265 388 297
rect 464 265 494 297
rect 548 265 578 297
rect 632 265 662 297
rect 716 265 746 297
rect 30 249 114 265
rect 30 215 40 249
rect 74 215 114 249
rect 30 199 114 215
rect 166 249 220 265
rect 166 215 176 249
rect 210 215 220 249
rect 166 199 220 215
rect 262 249 316 265
rect 262 215 272 249
rect 306 215 316 249
rect 262 199 316 215
rect 358 249 412 265
rect 358 215 368 249
rect 402 215 412 249
rect 358 199 412 215
rect 464 249 746 265
rect 464 215 474 249
rect 508 215 542 249
rect 576 215 610 249
rect 644 215 678 249
rect 712 215 746 249
rect 464 199 746 215
rect 84 177 114 199
rect 190 177 220 199
rect 274 177 304 199
rect 358 177 388 199
rect 464 177 494 199
rect 548 177 578 199
rect 632 177 662 199
rect 716 177 746 199
rect 84 21 114 47
rect 190 21 220 47
rect 274 21 304 47
rect 358 21 388 47
rect 464 21 494 47
rect 548 21 578 47
rect 632 21 662 47
rect 716 21 746 47
<< polycont >>
rect 40 215 74 249
rect 176 215 210 249
rect 272 215 306 249
rect 368 215 402 249
rect 474 215 508 249
rect 542 215 576 249
rect 610 215 644 249
rect 678 215 712 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 23 485 90 490
rect 23 451 40 485
rect 74 451 90 485
rect 401 477 451 527
rect 23 417 90 451
rect 23 383 40 417
rect 74 383 90 417
rect 23 349 90 383
rect 23 315 40 349
rect 74 333 90 349
rect 74 315 142 333
rect 23 299 142 315
rect 17 249 74 265
rect 17 215 40 249
rect 17 151 74 215
rect 108 165 142 299
rect 176 324 246 475
rect 280 357 344 475
rect 401 443 409 477
rect 443 443 451 477
rect 401 409 451 443
rect 401 375 409 409
rect 443 375 451 409
rect 401 359 451 375
rect 496 477 546 493
rect 496 443 504 477
rect 538 443 546 477
rect 496 409 546 443
rect 496 375 504 409
rect 538 375 546 409
rect 176 249 210 324
rect 280 290 322 357
rect 496 341 546 375
rect 580 477 630 527
rect 580 443 588 477
rect 622 443 630 477
rect 580 409 630 443
rect 580 375 588 409
rect 622 375 630 409
rect 580 359 630 375
rect 664 477 714 493
rect 664 443 672 477
rect 706 443 714 477
rect 664 409 714 443
rect 664 375 672 409
rect 706 375 714 409
rect 176 199 210 215
rect 256 249 322 290
rect 256 215 272 249
rect 306 215 322 249
rect 256 199 322 215
rect 368 289 455 323
rect 496 307 504 341
rect 538 325 546 341
rect 664 341 714 375
rect 748 477 798 527
rect 748 443 756 477
rect 790 443 798 477
rect 748 409 798 443
rect 748 375 756 409
rect 790 375 798 409
rect 748 359 798 375
rect 664 325 672 341
rect 538 307 672 325
rect 706 325 714 341
rect 706 307 811 325
rect 496 291 811 307
rect 368 249 402 289
rect 368 199 402 215
rect 436 215 474 249
rect 508 215 542 249
rect 576 215 610 249
rect 644 215 678 249
rect 712 215 728 249
rect 436 165 470 215
rect 762 181 811 291
rect 108 131 470 165
rect 504 163 811 181
rect 504 145 672 163
rect 24 101 74 117
rect 24 67 40 101
rect 24 17 74 67
rect 140 115 174 131
rect 314 115 348 131
rect 140 61 174 81
rect 214 63 230 97
rect 264 63 280 97
rect 214 17 280 63
rect 504 114 554 145
rect 314 61 348 81
rect 392 63 418 97
rect 452 63 468 97
rect 392 17 468 63
rect 538 80 554 114
rect 656 129 672 145
rect 706 145 811 163
rect 706 129 722 145
rect 504 51 554 80
rect 588 95 622 111
rect 588 17 622 61
rect 656 95 722 129
rect 656 61 672 95
rect 706 61 722 95
rect 656 51 722 61
rect 756 95 790 111
rect 756 17 790 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 304 425 338 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 304 357 338 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 212 357 246 391 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 396 289 430 323 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 212 425 246 459 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 28 221 62 255 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 764 153 798 187 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 or4_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1068202
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1060956
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.140 0.000 
<< end >>
