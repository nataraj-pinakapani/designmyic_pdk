magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 30 980 3247 1086
<< pwell >>
rect 15 10 3251 96
<< mvpsubdiff >>
rect 41 36 107 70
rect 141 36 175 70
rect 209 36 243 70
rect 277 36 311 70
rect 345 36 379 70
rect 413 36 447 70
rect 481 36 515 70
rect 549 36 583 70
rect 617 36 651 70
rect 685 36 719 70
rect 753 36 787 70
rect 821 36 855 70
rect 889 36 923 70
rect 957 36 991 70
rect 1025 36 1059 70
rect 1093 36 1127 70
rect 1161 36 1195 70
rect 1229 36 1263 70
rect 1297 36 1331 70
rect 1365 36 1399 70
rect 1433 36 1467 70
rect 1501 36 1535 70
rect 1569 36 1603 70
rect 1637 36 1671 70
rect 1705 36 1739 70
rect 1773 36 1807 70
rect 1841 36 1875 70
rect 1909 36 1943 70
rect 1977 36 2011 70
rect 2045 36 2079 70
rect 2113 36 2147 70
rect 2181 36 2215 70
rect 2249 36 2283 70
rect 2317 36 2351 70
rect 2385 36 2419 70
rect 2453 36 2487 70
rect 2521 36 2555 70
rect 2589 36 2623 70
rect 2657 36 2691 70
rect 2725 36 2759 70
rect 2793 36 2827 70
rect 2861 36 2895 70
rect 2929 36 2963 70
rect 2997 36 3031 70
rect 3065 36 3099 70
rect 3133 36 3167 70
rect 3201 36 3225 70
<< mvnsubdiff >>
rect 66 1016 93 1050
rect 127 1016 161 1050
rect 195 1016 229 1050
rect 263 1016 297 1050
rect 331 1016 365 1050
rect 399 1016 433 1050
rect 467 1016 501 1050
rect 535 1016 569 1050
rect 603 1016 637 1050
rect 671 1016 705 1050
rect 739 1016 773 1050
rect 807 1016 841 1050
rect 875 1016 909 1050
rect 943 1016 977 1050
rect 1011 1016 1045 1050
rect 1079 1016 1113 1050
rect 1147 1016 1181 1050
rect 1215 1016 1249 1050
rect 1283 1016 1317 1050
rect 1351 1016 1385 1050
rect 1419 1016 1453 1050
rect 1487 1016 1521 1050
rect 1555 1016 1589 1050
rect 1623 1016 1657 1050
rect 1691 1016 1725 1050
rect 1759 1016 1793 1050
rect 1827 1016 1861 1050
rect 1895 1016 1929 1050
rect 1963 1016 1997 1050
rect 2031 1016 2065 1050
rect 2099 1016 2133 1050
rect 2167 1016 2201 1050
rect 2235 1016 2269 1050
rect 2303 1016 2337 1050
rect 2371 1016 2405 1050
rect 2439 1016 2473 1050
rect 2507 1016 2541 1050
rect 2575 1016 2609 1050
rect 2643 1016 2677 1050
rect 2711 1016 2745 1050
rect 2779 1016 2813 1050
rect 2847 1016 2881 1050
rect 2915 1016 2949 1050
rect 2983 1016 3017 1050
rect 3051 1016 3085 1050
rect 3119 1016 3153 1050
rect 3187 1016 3211 1050
<< mvpsubdiffcont >>
rect 107 36 141 70
rect 175 36 209 70
rect 243 36 277 70
rect 311 36 345 70
rect 379 36 413 70
rect 447 36 481 70
rect 515 36 549 70
rect 583 36 617 70
rect 651 36 685 70
rect 719 36 753 70
rect 787 36 821 70
rect 855 36 889 70
rect 923 36 957 70
rect 991 36 1025 70
rect 1059 36 1093 70
rect 1127 36 1161 70
rect 1195 36 1229 70
rect 1263 36 1297 70
rect 1331 36 1365 70
rect 1399 36 1433 70
rect 1467 36 1501 70
rect 1535 36 1569 70
rect 1603 36 1637 70
rect 1671 36 1705 70
rect 1739 36 1773 70
rect 1807 36 1841 70
rect 1875 36 1909 70
rect 1943 36 1977 70
rect 2011 36 2045 70
rect 2079 36 2113 70
rect 2147 36 2181 70
rect 2215 36 2249 70
rect 2283 36 2317 70
rect 2351 36 2385 70
rect 2419 36 2453 70
rect 2487 36 2521 70
rect 2555 36 2589 70
rect 2623 36 2657 70
rect 2691 36 2725 70
rect 2759 36 2793 70
rect 2827 36 2861 70
rect 2895 36 2929 70
rect 2963 36 2997 70
rect 3031 36 3065 70
rect 3099 36 3133 70
rect 3167 36 3201 70
<< mvnsubdiffcont >>
rect 93 1016 127 1050
rect 161 1016 195 1050
rect 229 1016 263 1050
rect 297 1016 331 1050
rect 365 1016 399 1050
rect 433 1016 467 1050
rect 501 1016 535 1050
rect 569 1016 603 1050
rect 637 1016 671 1050
rect 705 1016 739 1050
rect 773 1016 807 1050
rect 841 1016 875 1050
rect 909 1016 943 1050
rect 977 1016 1011 1050
rect 1045 1016 1079 1050
rect 1113 1016 1147 1050
rect 1181 1016 1215 1050
rect 1249 1016 1283 1050
rect 1317 1016 1351 1050
rect 1385 1016 1419 1050
rect 1453 1016 1487 1050
rect 1521 1016 1555 1050
rect 1589 1016 1623 1050
rect 1657 1016 1691 1050
rect 1725 1016 1759 1050
rect 1793 1016 1827 1050
rect 1861 1016 1895 1050
rect 1929 1016 1963 1050
rect 1997 1016 2031 1050
rect 2065 1016 2099 1050
rect 2133 1016 2167 1050
rect 2201 1016 2235 1050
rect 2269 1016 2303 1050
rect 2337 1016 2371 1050
rect 2405 1016 2439 1050
rect 2473 1016 2507 1050
rect 2541 1016 2575 1050
rect 2609 1016 2643 1050
rect 2677 1016 2711 1050
rect 2745 1016 2779 1050
rect 2813 1016 2847 1050
rect 2881 1016 2915 1050
rect 2949 1016 2983 1050
rect 3017 1016 3051 1050
rect 3085 1016 3119 1050
rect 3153 1016 3187 1050
<< locali >>
rect 66 1016 93 1050
rect 127 1016 141 1050
rect 195 1016 213 1050
rect 263 1016 285 1050
rect 331 1016 357 1050
rect 399 1016 429 1050
rect 467 1016 501 1050
rect 535 1016 569 1050
rect 607 1016 637 1050
rect 679 1016 705 1050
rect 751 1016 773 1050
rect 823 1016 841 1050
rect 895 1016 909 1050
rect 967 1016 977 1050
rect 1039 1016 1045 1050
rect 1111 1016 1113 1050
rect 1147 1016 1149 1050
rect 1215 1016 1221 1050
rect 1283 1016 1293 1050
rect 1351 1016 1365 1050
rect 1419 1016 1437 1050
rect 1487 1016 1509 1050
rect 1555 1016 1581 1050
rect 1623 1016 1653 1050
rect 1691 1016 1725 1050
rect 1759 1016 1793 1050
rect 1831 1016 1861 1050
rect 1903 1016 1929 1050
rect 1975 1016 1997 1050
rect 2047 1016 2065 1050
rect 2119 1016 2133 1050
rect 2191 1016 2201 1050
rect 2263 1016 2269 1050
rect 2335 1016 2337 1050
rect 2371 1016 2373 1050
rect 2439 1016 2445 1050
rect 2507 1016 2517 1050
rect 2575 1016 2589 1050
rect 2643 1016 2661 1050
rect 2711 1016 2733 1050
rect 2779 1016 2805 1050
rect 2847 1016 2877 1050
rect 2915 1016 2949 1050
rect 2983 1016 3017 1050
rect 3055 1016 3085 1050
rect 3127 1016 3153 1050
rect 3199 1016 3211 1050
rect 3170 791 3208 825
rect 1248 747 1314 752
rect 888 721 922 726
rect 888 649 922 687
rect 536 628 570 633
rect 1248 713 1262 747
rect 1296 713 1314 747
rect 1248 675 1314 713
rect 1248 641 1262 675
rect 1296 641 1314 675
rect 250 563 284 568
rect 250 491 284 529
rect 536 556 570 594
rect 320 390 392 434
rect 623 430 657 435
rect 1248 434 1314 641
rect 1350 683 1384 688
rect 1350 611 1384 649
rect 1702 655 1736 660
rect 1702 583 1736 621
rect 2789 484 2827 518
rect 1609 464 1643 469
rect 127 356 165 390
rect 199 356 204 390
rect 320 356 331 390
rect 365 356 403 390
rect 437 356 446 390
rect 623 358 657 396
rect 958 390 1079 434
rect 1609 392 1643 430
rect 320 332 392 356
rect 765 356 803 390
rect 837 356 842 390
rect 958 356 968 390
rect 1002 356 1040 390
rect 1074 356 1079 390
rect 1465 356 1503 390
rect 1537 356 1542 390
rect 1702 435 1736 440
rect 1702 363 1736 401
rect 1915 398 1949 436
rect 2002 398 2036 436
rect 3069 463 3081 497
rect 3115 463 3135 497
rect 2138 401 2179 434
rect 2213 401 2254 434
rect 958 332 1079 356
rect 2138 363 2254 401
rect 2138 332 2179 363
rect 2213 332 2254 363
rect 2445 363 2479 401
rect 2531 401 2619 434
rect 2653 401 2780 434
rect 2531 363 2780 401
rect 2531 329 2619 363
rect 2653 329 2780 363
rect 3069 434 3135 463
rect 2899 363 2933 401
rect 3081 425 3115 434
rect 2531 322 2780 329
rect 2531 151 2607 322
rect 41 36 83 70
rect 141 36 155 70
rect 209 36 227 70
rect 277 36 299 70
rect 345 36 371 70
rect 413 36 443 70
rect 481 36 515 70
rect 549 36 583 70
rect 621 36 651 70
rect 693 36 719 70
rect 765 36 787 70
rect 837 36 855 70
rect 909 36 923 70
rect 981 36 991 70
rect 1053 36 1059 70
rect 1125 36 1127 70
rect 1161 36 1163 70
rect 1229 36 1235 70
rect 1297 36 1307 70
rect 1365 36 1379 70
rect 1433 36 1451 70
rect 1501 36 1523 70
rect 1569 36 1595 70
rect 1637 36 1667 70
rect 1705 36 1739 70
rect 1773 36 1807 70
rect 1845 36 1875 70
rect 1917 36 1943 70
rect 1989 36 2011 70
rect 2061 36 2079 70
rect 2133 36 2147 70
rect 2205 36 2215 70
rect 2277 36 2283 70
rect 2349 36 2351 70
rect 2385 36 2387 70
rect 2453 36 2459 70
rect 2521 36 2531 70
rect 2589 36 2603 70
rect 2657 36 2675 70
rect 2725 36 2747 70
rect 2793 36 2819 70
rect 2861 36 2891 70
rect 2929 36 2963 70
rect 2997 36 3031 70
rect 3069 36 3099 70
rect 3141 36 3167 70
rect 3213 36 3225 70
<< viali >>
rect 141 1016 161 1050
rect 161 1016 175 1050
rect 213 1016 229 1050
rect 229 1016 247 1050
rect 285 1016 297 1050
rect 297 1016 319 1050
rect 357 1016 365 1050
rect 365 1016 391 1050
rect 429 1016 433 1050
rect 433 1016 463 1050
rect 501 1016 535 1050
rect 573 1016 603 1050
rect 603 1016 607 1050
rect 645 1016 671 1050
rect 671 1016 679 1050
rect 717 1016 739 1050
rect 739 1016 751 1050
rect 789 1016 807 1050
rect 807 1016 823 1050
rect 861 1016 875 1050
rect 875 1016 895 1050
rect 933 1016 943 1050
rect 943 1016 967 1050
rect 1005 1016 1011 1050
rect 1011 1016 1039 1050
rect 1077 1016 1079 1050
rect 1079 1016 1111 1050
rect 1149 1016 1181 1050
rect 1181 1016 1183 1050
rect 1221 1016 1249 1050
rect 1249 1016 1255 1050
rect 1293 1016 1317 1050
rect 1317 1016 1327 1050
rect 1365 1016 1385 1050
rect 1385 1016 1399 1050
rect 1437 1016 1453 1050
rect 1453 1016 1471 1050
rect 1509 1016 1521 1050
rect 1521 1016 1543 1050
rect 1581 1016 1589 1050
rect 1589 1016 1615 1050
rect 1653 1016 1657 1050
rect 1657 1016 1687 1050
rect 1725 1016 1759 1050
rect 1797 1016 1827 1050
rect 1827 1016 1831 1050
rect 1869 1016 1895 1050
rect 1895 1016 1903 1050
rect 1941 1016 1963 1050
rect 1963 1016 1975 1050
rect 2013 1016 2031 1050
rect 2031 1016 2047 1050
rect 2085 1016 2099 1050
rect 2099 1016 2119 1050
rect 2157 1016 2167 1050
rect 2167 1016 2191 1050
rect 2229 1016 2235 1050
rect 2235 1016 2263 1050
rect 2301 1016 2303 1050
rect 2303 1016 2335 1050
rect 2373 1016 2405 1050
rect 2405 1016 2407 1050
rect 2445 1016 2473 1050
rect 2473 1016 2479 1050
rect 2517 1016 2541 1050
rect 2541 1016 2551 1050
rect 2589 1016 2609 1050
rect 2609 1016 2623 1050
rect 2661 1016 2677 1050
rect 2677 1016 2695 1050
rect 2733 1016 2745 1050
rect 2745 1016 2767 1050
rect 2805 1016 2813 1050
rect 2813 1016 2839 1050
rect 2877 1016 2881 1050
rect 2881 1016 2911 1050
rect 2949 1016 2983 1050
rect 3021 1016 3051 1050
rect 3051 1016 3055 1050
rect 3093 1016 3119 1050
rect 3119 1016 3127 1050
rect 3165 1016 3187 1050
rect 3187 1016 3199 1050
rect 3136 791 3170 825
rect 3208 791 3242 825
rect 888 687 922 721
rect 536 594 570 628
rect 888 615 922 649
rect 1262 713 1296 747
rect 1262 641 1296 675
rect 250 529 284 563
rect 536 522 570 556
rect 250 457 284 491
rect 1350 649 1384 683
rect 1350 577 1384 611
rect 1702 621 1736 655
rect 1702 549 1736 583
rect 2755 484 2789 518
rect 2827 484 2861 518
rect 623 396 657 430
rect 93 356 127 390
rect 165 356 199 390
rect 331 356 365 390
rect 403 356 437 390
rect 1609 430 1643 464
rect 623 324 657 358
rect 731 356 765 390
rect 803 356 837 390
rect 968 356 1002 390
rect 1040 356 1074 390
rect 1431 356 1465 390
rect 1503 356 1537 390
rect 1609 358 1643 392
rect 1702 401 1736 435
rect 1915 436 1949 470
rect 1915 364 1949 398
rect 2002 436 2036 470
rect 3081 463 3115 497
rect 2002 364 2036 398
rect 2179 401 2213 435
rect 1702 329 1736 363
rect 2179 329 2213 363
rect 2445 401 2479 435
rect 2445 329 2479 363
rect 2619 401 2653 435
rect 2619 329 2653 363
rect 2899 401 2933 435
rect 3081 391 3115 425
rect 2899 329 2933 363
rect 83 36 107 70
rect 107 36 117 70
rect 155 36 175 70
rect 175 36 189 70
rect 227 36 243 70
rect 243 36 261 70
rect 299 36 311 70
rect 311 36 333 70
rect 371 36 379 70
rect 379 36 405 70
rect 443 36 447 70
rect 447 36 477 70
rect 515 36 549 70
rect 587 36 617 70
rect 617 36 621 70
rect 659 36 685 70
rect 685 36 693 70
rect 731 36 753 70
rect 753 36 765 70
rect 803 36 821 70
rect 821 36 837 70
rect 875 36 889 70
rect 889 36 909 70
rect 947 36 957 70
rect 957 36 981 70
rect 1019 36 1025 70
rect 1025 36 1053 70
rect 1091 36 1093 70
rect 1093 36 1125 70
rect 1163 36 1195 70
rect 1195 36 1197 70
rect 1235 36 1263 70
rect 1263 36 1269 70
rect 1307 36 1331 70
rect 1331 36 1341 70
rect 1379 36 1399 70
rect 1399 36 1413 70
rect 1451 36 1467 70
rect 1467 36 1485 70
rect 1523 36 1535 70
rect 1535 36 1557 70
rect 1595 36 1603 70
rect 1603 36 1629 70
rect 1667 36 1671 70
rect 1671 36 1701 70
rect 1739 36 1773 70
rect 1811 36 1841 70
rect 1841 36 1845 70
rect 1883 36 1909 70
rect 1909 36 1917 70
rect 1955 36 1977 70
rect 1977 36 1989 70
rect 2027 36 2045 70
rect 2045 36 2061 70
rect 2099 36 2113 70
rect 2113 36 2133 70
rect 2171 36 2181 70
rect 2181 36 2205 70
rect 2243 36 2249 70
rect 2249 36 2277 70
rect 2315 36 2317 70
rect 2317 36 2349 70
rect 2387 36 2419 70
rect 2419 36 2421 70
rect 2459 36 2487 70
rect 2487 36 2493 70
rect 2531 36 2555 70
rect 2555 36 2565 70
rect 2603 36 2623 70
rect 2623 36 2637 70
rect 2675 36 2691 70
rect 2691 36 2709 70
rect 2747 36 2759 70
rect 2759 36 2781 70
rect 2819 36 2827 70
rect 2827 36 2853 70
rect 2891 36 2895 70
rect 2895 36 2925 70
rect 2963 36 2997 70
rect 3035 36 3065 70
rect 3065 36 3069 70
rect 3107 36 3133 70
rect 3133 36 3141 70
rect 3179 36 3201 70
rect 3201 36 3213 70
<< metal1 >>
rect 66 1050 3211 1062
rect 66 1016 141 1050
rect 175 1016 213 1050
rect 247 1016 285 1050
rect 319 1016 357 1050
rect 391 1016 429 1050
rect 463 1016 501 1050
rect 535 1016 573 1050
rect 607 1016 645 1050
rect 679 1016 717 1050
rect 751 1016 789 1050
rect 823 1016 861 1050
rect 895 1016 933 1050
rect 967 1016 1005 1050
rect 1039 1016 1077 1050
rect 1111 1016 1149 1050
rect 1183 1016 1221 1050
rect 1255 1016 1293 1050
rect 1327 1016 1365 1050
rect 1399 1016 1437 1050
rect 1471 1016 1509 1050
rect 1543 1016 1581 1050
rect 1615 1016 1653 1050
rect 1687 1016 1725 1050
rect 1759 1016 1797 1050
rect 1831 1016 1869 1050
rect 1903 1016 1941 1050
rect 1975 1016 2013 1050
rect 2047 1016 2085 1050
rect 2119 1016 2157 1050
rect 2191 1016 2229 1050
rect 2263 1016 2301 1050
rect 2335 1016 2373 1050
rect 2407 1016 2445 1050
rect 2479 1016 2517 1050
rect 2551 1016 2589 1050
rect 2623 1016 2661 1050
rect 2695 1016 2733 1050
rect 2767 1016 2805 1050
rect 2839 1016 2877 1050
rect 2911 1016 2949 1050
rect 2983 1016 3021 1050
rect 3055 1016 3093 1050
rect 3127 1016 3165 1050
rect 3199 1016 3211 1050
rect 66 1004 3211 1016
rect 245 859 2632 1004
rect 3124 825 3254 831
rect 3124 791 3136 825
rect 3170 791 3208 825
rect 3242 791 3254 825
rect 3124 785 3254 791
rect 1256 747 1302 764
rect 882 721 928 738
rect 882 687 888 721
rect 922 687 928 721
rect 882 675 928 687
rect 1256 713 1262 747
rect 1296 713 1302 747
tri 928 675 936 683 sw
rect 1256 675 1302 713
rect 882 649 936 675
tri 936 649 962 675 sw
rect 530 628 576 645
rect 530 594 536 628
rect 570 594 576 628
rect 882 615 888 649
rect 922 641 1178 649
tri 1178 641 1186 649 sw
rect 1256 641 1262 675
rect 1296 641 1302 675
rect 922 629 1186 641
tri 1186 629 1198 641 sw
rect 1256 629 1302 641
rect 1344 683 1390 700
rect 1344 649 1350 683
rect 1384 649 1390 683
rect 922 621 1198 629
tri 1198 621 1206 629 sw
rect 922 615 1206 621
rect 882 611 1206 615
tri 1206 611 1216 621 sw
rect 1344 617 1390 649
rect 1696 655 1742 672
rect 1696 621 1702 655
rect 1736 621 1742 655
tri 1390 617 1393 620 sw
rect 1344 611 1393 617
rect 882 603 1216 611
tri 1216 603 1224 611 sw
rect 244 563 290 580
rect 244 529 250 563
rect 284 529 290 563
rect 244 522 290 529
rect 530 577 576 594
tri 1158 590 1171 603 ne
rect 1171 590 1224 603
tri 1224 590 1237 603 sw
tri 576 577 589 590 sw
tri 1171 583 1178 590 ne
rect 1178 583 1237 590
tri 1237 583 1244 590 sw
tri 1178 577 1184 583 ne
rect 1184 577 1244 583
tri 1244 577 1250 583 sw
rect 1344 577 1350 611
rect 1384 583 1393 611
tri 1393 583 1427 617 sw
rect 1696 583 1742 621
rect 1384 577 1427 583
rect 530 565 589 577
tri 589 565 601 577 sw
tri 1184 565 1196 577 ne
rect 1196 565 1250 577
tri 1250 565 1262 577 sw
rect 1344 565 1427 577
rect 530 556 601 565
tri 601 556 610 565 sw
tri 1196 556 1205 565 ne
rect 1205 556 1262 565
tri 1262 556 1271 565 sw
tri 1377 556 1386 565 ne
rect 1386 556 1427 565
tri 290 522 293 525 sw
rect 530 522 536 556
rect 570 555 815 556
tri 815 555 816 556 sw
tri 1205 555 1206 556 ne
rect 1206 555 1271 556
tri 1271 555 1272 556 sw
tri 1386 555 1387 556 ne
rect 1387 555 1427 556
rect 570 554 816 555
tri 816 554 817 555 sw
tri 1206 554 1207 555 ne
rect 1207 554 1272 555
tri 1272 554 1273 555 sw
tri 1387 554 1388 555 ne
rect 1388 554 1427 555
rect 570 553 817 554
tri 817 553 818 554 sw
tri 1207 553 1208 554 ne
rect 1208 553 1273 554
tri 1273 553 1274 554 sw
tri 1388 553 1389 554 ne
rect 1389 553 1427 554
rect 570 552 818 553
tri 818 552 819 553 sw
tri 1208 552 1209 553 ne
rect 1209 552 1274 553
tri 1274 552 1275 553 sw
tri 1389 552 1390 553 ne
rect 1390 552 1427 553
rect 570 551 819 552
tri 819 551 820 552 sw
tri 1209 551 1210 552 ne
rect 1210 551 1275 552
tri 1275 551 1276 552 sw
tri 1390 551 1391 552 ne
rect 1391 551 1427 552
rect 570 550 820 551
tri 820 550 821 551 sw
tri 1210 550 1211 551 ne
rect 1211 550 1276 551
tri 1276 550 1277 551 sw
tri 1391 550 1392 551 ne
rect 1392 550 1427 551
rect 570 549 821 550
tri 821 549 822 550 sw
tri 1211 549 1212 550 ne
rect 1212 549 1277 550
tri 1277 549 1278 550 sw
tri 1392 549 1393 550 ne
rect 1393 549 1427 550
tri 1427 549 1461 583 sw
rect 1696 549 1702 583
rect 1736 549 1742 583
rect 570 548 822 549
tri 822 548 823 549 sw
tri 1212 548 1213 549 ne
rect 1213 548 1278 549
tri 1278 548 1279 549 sw
tri 1393 548 1394 549 ne
rect 1394 548 1461 549
rect 570 547 823 548
tri 823 547 824 548 sw
tri 1213 547 1214 548 ne
rect 1214 547 1279 548
tri 1279 547 1280 548 sw
tri 1394 547 1395 548 ne
rect 1395 547 1461 548
rect 570 546 824 547
tri 824 546 825 547 sw
tri 1214 546 1215 547 ne
rect 1215 546 1280 547
tri 1280 546 1281 547 sw
tri 1395 546 1396 547 ne
rect 1396 546 1461 547
rect 570 545 825 546
tri 825 545 826 546 sw
tri 1215 545 1216 546 ne
rect 1216 545 1281 546
tri 1281 545 1282 546 sw
tri 1396 545 1397 546 ne
rect 1397 545 1461 546
rect 570 544 826 545
tri 826 544 827 545 sw
tri 1216 544 1217 545 ne
rect 1217 544 1282 545
tri 1282 544 1283 545 sw
tri 1397 544 1398 545 ne
rect 1398 544 1461 545
rect 570 543 827 544
tri 827 543 828 544 sw
tri 1217 543 1218 544 ne
rect 1218 543 1283 544
tri 1283 543 1284 544 sw
tri 1398 543 1399 544 ne
rect 1399 543 1461 544
rect 570 542 828 543
tri 828 542 829 543 sw
tri 1218 542 1219 543 ne
rect 1219 542 1284 543
tri 1284 542 1285 543 sw
tri 1399 542 1400 543 ne
rect 1400 542 1461 543
rect 570 541 829 542
tri 829 541 830 542 sw
tri 1219 541 1220 542 ne
rect 1220 541 1285 542
tri 1285 541 1286 542 sw
tri 1400 541 1401 542 ne
rect 1401 541 1461 542
rect 570 540 830 541
tri 830 540 831 541 sw
tri 1220 540 1221 541 ne
rect 1221 540 1286 541
tri 1286 540 1287 541 sw
tri 1401 540 1402 541 ne
rect 1402 540 1461 541
rect 570 539 831 540
tri 831 539 832 540 sw
tri 1221 539 1222 540 ne
rect 1222 539 1287 540
tri 1287 539 1288 540 sw
tri 1402 539 1403 540 ne
rect 1403 539 1461 540
rect 570 538 832 539
tri 832 538 833 539 sw
tri 1222 538 1223 539 ne
rect 1223 538 1288 539
tri 1288 538 1289 539 sw
tri 1403 538 1404 539 ne
rect 1404 538 1461 539
rect 570 537 833 538
tri 833 537 834 538 sw
tri 1223 537 1224 538 ne
rect 1224 537 1289 538
tri 1289 537 1290 538 sw
tri 1404 537 1405 538 ne
rect 1405 537 1461 538
rect 570 536 834 537
tri 834 536 835 537 sw
tri 1224 536 1225 537 ne
rect 1225 536 1290 537
tri 1290 536 1291 537 sw
tri 1405 536 1406 537 ne
rect 1406 536 1461 537
rect 570 535 835 536
tri 835 535 836 536 sw
tri 1225 535 1226 536 ne
rect 1226 535 1291 536
tri 1291 535 1292 536 sw
tri 1406 535 1407 536 ne
rect 1407 535 1461 536
rect 570 534 836 535
tri 836 534 837 535 sw
tri 1226 534 1227 535 ne
rect 1227 534 1292 535
tri 1292 534 1293 535 sw
tri 1407 534 1408 535 ne
rect 1408 534 1461 535
rect 570 533 837 534
tri 837 533 838 534 sw
tri 1227 533 1228 534 ne
rect 1228 533 1293 534
tri 1293 533 1294 534 sw
tri 1408 533 1409 534 ne
rect 1409 533 1461 534
rect 570 532 838 533
tri 838 532 839 533 sw
tri 1228 532 1229 533 ne
rect 1229 532 1294 533
tri 1294 532 1295 533 sw
tri 1409 532 1410 533 ne
rect 1410 532 1461 533
rect 570 531 839 532
tri 839 531 840 532 sw
tri 1229 531 1230 532 ne
rect 1230 531 1295 532
tri 1295 531 1296 532 sw
tri 1410 531 1411 532 ne
rect 1411 531 1461 532
rect 570 530 840 531
tri 840 530 841 531 sw
tri 1230 530 1231 531 ne
rect 1231 530 1296 531
tri 1296 530 1297 531 sw
tri 1411 530 1412 531 ne
rect 1412 530 1461 531
rect 570 529 841 530
tri 841 529 842 530 sw
tri 1231 529 1232 530 ne
rect 1232 529 1297 530
tri 1297 529 1298 530 sw
tri 1412 529 1413 530 ne
rect 1413 529 1461 530
rect 570 528 842 529
tri 842 528 843 529 sw
tri 1232 528 1233 529 ne
rect 1233 528 1298 529
tri 1298 528 1299 529 sw
tri 1413 528 1414 529 ne
rect 1414 528 1461 529
rect 570 527 843 528
tri 843 527 844 528 sw
tri 1233 527 1234 528 ne
rect 1234 527 1299 528
tri 1299 527 1300 528 sw
tri 1414 527 1415 528 ne
rect 1415 527 1461 528
rect 570 526 844 527
tri 844 526 845 527 sw
tri 1234 526 1235 527 ne
rect 1235 526 1300 527
tri 1300 526 1301 527 sw
tri 1415 526 1416 527 ne
rect 1416 526 1461 527
rect 570 525 845 526
tri 845 525 846 526 sw
tri 1235 525 1236 526 ne
rect 1236 525 1301 526
tri 1301 525 1302 526 sw
tri 1416 525 1417 526 ne
rect 1417 525 1461 526
rect 570 524 846 525
tri 846 524 847 525 sw
tri 1236 524 1237 525 ne
rect 1237 524 1302 525
tri 1302 524 1303 525 sw
tri 1417 524 1418 525 ne
rect 1418 524 1461 525
rect 570 523 847 524
tri 847 523 848 524 sw
tri 1237 523 1238 524 ne
rect 1238 523 1303 524
tri 1303 523 1304 524 sw
tri 1418 523 1419 524 ne
rect 1419 523 1461 524
rect 570 522 848 523
tri 848 522 849 523 sw
tri 1238 522 1239 523 ne
rect 1239 522 1304 523
tri 1304 522 1305 523 sw
tri 1419 522 1420 523 ne
rect 1420 522 1461 523
rect 244 518 293 522
tri 293 518 297 522 sw
rect 530 521 849 522
tri 849 521 850 522 sw
tri 1239 521 1240 522 ne
rect 1240 521 1305 522
tri 1305 521 1306 522 sw
tri 1420 521 1421 522 ne
rect 1421 521 1461 522
rect 530 520 850 521
tri 850 520 851 521 sw
tri 1240 520 1241 521 ne
rect 1241 520 1306 521
tri 1306 520 1307 521 sw
tri 1421 520 1422 521 ne
rect 1422 520 1461 521
rect 530 519 851 520
tri 851 519 852 520 sw
tri 1241 519 1242 520 ne
rect 1242 519 1307 520
tri 1307 519 1308 520 sw
tri 1422 519 1423 520 ne
rect 1423 519 1461 520
rect 530 518 852 519
tri 852 518 853 519 sw
tri 1242 518 1243 519 ne
rect 1243 518 1308 519
tri 1308 518 1309 519 sw
tri 1423 518 1424 519 ne
rect 1424 518 1461 519
tri 1461 518 1492 549 sw
rect 1696 537 1742 549
tri 3065 524 3069 528 se
rect 2743 518 3121 524
rect 244 510 297 518
tri 297 510 305 518 sw
rect 530 517 853 518
tri 853 517 854 518 sw
tri 1243 517 1244 518 ne
rect 1244 517 1309 518
tri 1309 517 1310 518 sw
tri 1424 517 1425 518 ne
rect 1425 517 1492 518
rect 530 516 854 517
tri 854 516 855 517 sw
tri 1244 516 1245 517 ne
rect 1245 516 1310 517
tri 1310 516 1311 517 sw
tri 1425 516 1426 517 ne
rect 1426 516 1492 517
rect 530 515 855 516
tri 855 515 856 516 sw
tri 1245 515 1246 516 ne
rect 1246 515 1311 516
tri 1311 515 1312 516 sw
tri 1426 515 1427 516 ne
rect 1427 515 1492 516
rect 530 514 856 515
tri 856 514 857 515 sw
tri 1246 514 1247 515 ne
rect 1247 514 1312 515
tri 1312 514 1313 515 sw
tri 1427 514 1428 515 ne
rect 1428 514 1492 515
rect 530 513 857 514
tri 857 513 858 514 sw
tri 1247 513 1248 514 ne
rect 1248 513 1313 514
tri 1313 513 1314 514 sw
tri 1428 513 1429 514 ne
rect 1429 513 1492 514
rect 530 512 858 513
tri 858 512 859 513 sw
tri 1248 512 1249 513 ne
rect 1249 512 1314 513
tri 1314 512 1315 513 sw
tri 1429 512 1430 513 ne
rect 1430 512 1492 513
rect 530 511 859 512
tri 859 511 860 512 sw
tri 1249 511 1250 512 ne
rect 1250 511 1315 512
tri 1315 511 1316 512 sw
tri 1430 511 1431 512 ne
rect 1431 511 1492 512
rect 530 510 860 511
tri 860 510 861 511 sw
tri 1250 510 1251 511 ne
rect 1251 510 1316 511
tri 1316 510 1317 511 sw
tri 1431 510 1432 511 ne
rect 1432 510 1492 511
rect 244 491 305 510
tri 305 491 324 510 sw
tri 795 509 796 510 ne
rect 796 509 861 510
tri 861 509 862 510 sw
tri 1251 509 1252 510 ne
rect 1252 509 1317 510
tri 1317 509 1318 510 sw
tri 1432 509 1433 510 ne
rect 1433 509 1492 510
tri 796 508 797 509 ne
rect 797 508 862 509
tri 862 508 863 509 sw
tri 1252 508 1253 509 ne
rect 1253 508 1318 509
tri 1318 508 1319 509 sw
tri 1433 508 1434 509 ne
rect 1434 508 1492 509
tri 797 507 798 508 ne
rect 798 507 863 508
tri 863 507 864 508 sw
tri 1253 507 1254 508 ne
rect 1254 507 1319 508
tri 1319 507 1320 508 sw
tri 1434 507 1435 508 ne
rect 1435 507 1492 508
tri 798 506 799 507 ne
rect 799 506 864 507
tri 864 506 865 507 sw
tri 1254 506 1255 507 ne
rect 1255 506 1320 507
tri 1320 506 1321 507 sw
tri 1435 506 1436 507 ne
rect 1436 506 1492 507
tri 799 505 800 506 ne
rect 800 505 865 506
tri 865 505 866 506 sw
tri 1255 505 1256 506 ne
rect 1256 505 1321 506
tri 1321 505 1322 506 sw
tri 1436 505 1437 506 ne
rect 1437 505 1492 506
tri 800 504 801 505 ne
rect 801 504 866 505
tri 866 504 867 505 sw
tri 1256 504 1257 505 ne
rect 1257 504 1322 505
tri 1322 504 1323 505 sw
tri 1437 504 1438 505 ne
rect 1438 504 1492 505
tri 801 503 802 504 ne
rect 802 503 867 504
tri 867 503 868 504 sw
tri 1257 503 1258 504 ne
rect 1258 503 1323 504
tri 1323 503 1324 504 sw
tri 1438 503 1439 504 ne
rect 1439 503 1492 504
tri 802 502 803 503 ne
rect 803 502 868 503
tri 868 502 869 503 sw
tri 1258 502 1259 503 ne
rect 1259 502 1324 503
tri 1324 502 1325 503 sw
tri 1439 502 1440 503 ne
rect 1440 502 1492 503
tri 803 501 804 502 ne
rect 804 501 869 502
tri 869 501 870 502 sw
tri 1259 501 1260 502 ne
rect 1260 501 1325 502
tri 1325 501 1326 502 sw
tri 1440 501 1441 502 ne
rect 1441 501 1492 502
tri 804 500 805 501 ne
rect 805 500 870 501
tri 870 500 871 501 sw
tri 1260 500 1261 501 ne
rect 1261 500 1326 501
tri 1326 500 1327 501 sw
tri 1441 500 1442 501 ne
rect 1442 500 1492 501
tri 805 499 806 500 ne
rect 806 499 871 500
tri 871 499 872 500 sw
tri 1261 499 1262 500 ne
rect 1262 499 1327 500
tri 1327 499 1328 500 sw
tri 1442 499 1443 500 ne
rect 1443 499 1492 500
tri 806 498 807 499 ne
rect 807 498 872 499
tri 872 498 873 499 sw
tri 1262 498 1263 499 ne
rect 1263 498 1328 499
tri 1328 498 1329 499 sw
tri 1443 498 1444 499 ne
rect 1444 498 1492 499
tri 807 497 808 498 ne
rect 808 497 873 498
tri 873 497 874 498 sw
tri 1263 497 1264 498 ne
rect 1264 497 1329 498
tri 1329 497 1330 498 sw
tri 1444 497 1445 498 ne
rect 1445 497 1492 498
tri 808 496 809 497 ne
rect 809 496 874 497
tri 874 496 875 497 sw
tri 1264 496 1265 497 ne
rect 1265 496 1330 497
tri 1330 496 1331 497 sw
tri 1445 496 1446 497 ne
rect 1446 496 1492 497
tri 809 495 810 496 ne
rect 810 495 875 496
tri 875 495 876 496 sw
tri 1265 495 1266 496 ne
rect 1266 495 1331 496
tri 1331 495 1332 496 sw
tri 1446 495 1447 496 ne
rect 1447 495 1492 496
tri 810 494 811 495 ne
rect 811 494 876 495
tri 876 494 877 495 sw
tri 1266 494 1267 495 ne
rect 1267 494 1332 495
tri 1332 494 1333 495 sw
tri 1447 494 1448 495 ne
rect 1448 494 1492 495
tri 811 493 812 494 ne
rect 812 493 877 494
tri 877 493 878 494 sw
tri 1267 493 1268 494 ne
rect 1268 493 1333 494
tri 1333 493 1334 494 sw
tri 1448 493 1449 494 ne
rect 1449 493 1492 494
tri 812 492 813 493 ne
rect 813 492 878 493
tri 878 492 879 493 sw
tri 1268 492 1269 493 ne
rect 1269 492 1334 493
tri 1334 492 1335 493 sw
tri 1449 492 1450 493 ne
rect 1450 492 1492 493
tri 813 491 814 492 ne
rect 814 491 879 492
tri 879 491 880 492 sw
tri 1269 491 1270 492 ne
rect 1270 491 1335 492
tri 1335 491 1336 492 sw
tri 1450 491 1451 492 ne
rect 1451 491 1492 492
rect 244 457 250 491
rect 284 490 478 491
tri 478 490 479 491 sw
tri 814 490 815 491 ne
rect 815 490 880 491
tri 880 490 881 491 sw
tri 1270 490 1271 491 ne
rect 1271 490 1336 491
tri 1336 490 1337 491 sw
tri 1451 490 1452 491 ne
rect 1452 490 1492 491
rect 284 484 479 490
tri 479 484 485 490 sw
tri 815 489 816 490 ne
rect 816 489 881 490
tri 881 489 882 490 sw
tri 1271 489 1272 490 ne
rect 1272 489 1337 490
tri 1337 489 1338 490 sw
tri 1452 489 1453 490 ne
rect 1453 489 1492 490
tri 816 488 817 489 ne
rect 817 488 882 489
tri 882 488 883 489 sw
tri 1272 488 1273 489 ne
rect 1273 488 1338 489
tri 1338 488 1339 489 sw
tri 1453 488 1454 489 ne
rect 1454 488 1492 489
tri 817 487 818 488 ne
rect 818 487 883 488
tri 883 487 884 488 sw
tri 1273 487 1274 488 ne
rect 1274 487 1339 488
tri 1339 487 1340 488 sw
tri 1454 487 1455 488 ne
rect 1455 487 1492 488
tri 818 486 819 487 ne
rect 819 486 884 487
tri 884 486 885 487 sw
tri 1274 486 1275 487 ne
rect 1275 486 1340 487
tri 1340 486 1341 487 sw
tri 1455 486 1456 487 ne
rect 1456 486 1492 487
tri 819 485 820 486 ne
rect 820 485 885 486
tri 885 485 886 486 sw
tri 1275 485 1276 486 ne
rect 1276 485 1341 486
tri 1341 485 1342 486 sw
tri 1456 485 1457 486 ne
rect 1457 485 1492 486
tri 820 484 821 485 ne
rect 821 484 886 485
tri 886 484 887 485 sw
tri 1276 484 1277 485 ne
rect 1277 484 1342 485
tri 1342 484 1343 485 sw
tri 1457 484 1458 485 ne
rect 1458 484 1492 485
tri 1492 484 1526 518 sw
rect 2743 484 2755 518
rect 2789 484 2827 518
rect 2861 497 3121 518
rect 2861 484 3081 497
rect 284 470 485 484
tri 485 470 499 484 sw
tri 821 483 822 484 ne
rect 822 483 887 484
tri 887 483 888 484 sw
tri 1277 483 1278 484 ne
rect 1278 483 1343 484
tri 1343 483 1344 484 sw
tri 1458 483 1459 484 ne
rect 1459 483 1526 484
tri 822 482 823 483 ne
rect 823 482 888 483
tri 888 482 889 483 sw
tri 1278 482 1279 483 ne
rect 1279 482 1344 483
tri 1344 482 1345 483 sw
tri 1459 482 1460 483 ne
rect 1460 482 1526 483
tri 823 481 824 482 ne
rect 824 481 889 482
tri 889 481 890 482 sw
tri 1279 481 1280 482 ne
rect 1280 481 1345 482
tri 1345 481 1346 482 sw
tri 1460 481 1461 482 ne
rect 1461 481 1526 482
tri 1526 481 1529 484 sw
tri 824 480 825 481 ne
rect 825 480 890 481
tri 890 480 891 481 sw
tri 1280 480 1281 481 ne
rect 1281 480 1346 481
tri 1346 480 1347 481 sw
tri 1461 480 1462 481 ne
rect 1462 480 1649 481
tri 825 479 826 480 ne
rect 826 479 891 480
tri 891 479 892 480 sw
tri 1281 479 1282 480 ne
rect 1282 479 1347 480
tri 1347 479 1348 480 sw
tri 1462 479 1463 480 ne
rect 1463 479 1649 480
tri 826 478 827 479 ne
rect 827 478 892 479
tri 892 478 893 479 sw
tri 1282 478 1283 479 ne
rect 1283 478 1348 479
tri 1348 478 1349 479 sw
tri 1463 478 1464 479 ne
rect 1464 478 1649 479
tri 827 477 828 478 ne
rect 828 477 893 478
tri 893 477 894 478 sw
tri 1283 477 1284 478 ne
rect 1284 477 1349 478
tri 1349 477 1350 478 sw
tri 1464 477 1465 478 ne
rect 1465 477 1649 478
tri 828 476 829 477 ne
rect 829 476 894 477
tri 894 476 895 477 sw
tri 1284 476 1285 477 ne
rect 1285 476 1350 477
tri 1350 476 1351 477 sw
tri 1465 476 1466 477 ne
rect 1466 476 1649 477
tri 829 475 830 476 ne
rect 830 475 895 476
tri 895 475 896 476 sw
tri 1285 475 1286 476 ne
rect 1286 475 1351 476
tri 1351 475 1352 476 sw
tri 1466 475 1467 476 ne
rect 1467 475 1649 476
tri 830 474 831 475 ne
rect 831 474 896 475
tri 896 474 897 475 sw
tri 1286 474 1287 475 ne
rect 1287 474 1352 475
tri 1352 474 1353 475 sw
tri 1467 474 1468 475 ne
rect 1468 474 1649 475
tri 831 473 832 474 ne
rect 832 473 897 474
tri 897 473 898 474 sw
tri 1287 473 1288 474 ne
rect 1288 473 1353 474
tri 1353 473 1354 474 sw
tri 1468 473 1469 474 ne
rect 1469 473 1649 474
tri 832 472 833 473 ne
rect 833 472 898 473
tri 898 472 899 473 sw
tri 1288 472 1289 473 ne
rect 1289 472 1354 473
tri 1354 472 1355 473 sw
tri 1469 472 1470 473 ne
rect 1470 472 1649 473
tri 833 471 834 472 ne
rect 834 471 899 472
tri 899 471 900 472 sw
tri 1289 471 1290 472 ne
rect 1290 471 1355 472
tri 1355 471 1356 472 sw
tri 1470 471 1471 472 ne
rect 1471 471 1649 472
tri 834 470 835 471 ne
rect 835 470 900 471
tri 900 470 901 471 sw
tri 1290 470 1291 471 ne
rect 1291 470 1356 471
tri 1356 470 1357 471 sw
tri 1471 470 1472 471 ne
rect 1472 470 1649 471
rect 284 464 499 470
tri 499 464 505 470 sw
tri 835 469 836 470 ne
rect 836 469 901 470
tri 901 469 902 470 sw
tri 1291 469 1292 470 ne
rect 1292 469 1357 470
tri 1357 469 1358 470 sw
tri 1472 469 1473 470 ne
rect 1473 469 1649 470
tri 836 468 837 469 ne
rect 837 468 902 469
tri 902 468 903 469 sw
tri 1292 468 1293 469 ne
rect 1293 468 1358 469
tri 1358 468 1359 469 sw
tri 1473 468 1474 469 ne
rect 1474 468 1649 469
tri 837 467 838 468 ne
rect 838 467 903 468
tri 903 467 904 468 sw
tri 1293 467 1294 468 ne
rect 1294 467 1359 468
tri 1359 467 1360 468 sw
tri 1474 467 1475 468 ne
rect 1475 467 1649 468
tri 838 466 839 467 ne
rect 839 466 904 467
tri 904 466 905 467 sw
tri 1294 466 1295 467 ne
rect 1295 466 1360 467
tri 1360 466 1361 467 sw
tri 1475 466 1476 467 ne
rect 1476 466 1649 467
tri 839 465 840 466 ne
rect 840 465 905 466
tri 905 465 906 466 sw
tri 1295 465 1296 466 ne
rect 1296 465 1361 466
tri 1361 465 1362 466 sw
tri 1476 465 1477 466 ne
rect 1477 465 1649 466
tri 840 464 841 465 ne
rect 841 464 906 465
tri 906 464 907 465 sw
tri 1296 464 1297 465 ne
rect 1297 464 1362 465
tri 1362 464 1363 465 sw
tri 1477 464 1478 465 ne
rect 1478 464 1649 465
rect 284 457 505 464
rect 244 447 505 457
tri 505 447 522 464 sw
tri 841 463 842 464 ne
rect 842 463 907 464
tri 907 463 908 464 sw
tri 1297 463 1298 464 ne
rect 1298 463 1363 464
tri 1363 463 1364 464 sw
tri 1478 463 1479 464 ne
rect 1479 463 1609 464
tri 842 462 843 463 ne
rect 843 462 908 463
tri 908 462 909 463 sw
tri 1298 462 1299 463 ne
rect 1299 462 1364 463
tri 1364 462 1365 463 sw
tri 1479 462 1480 463 ne
rect 1480 462 1609 463
tri 843 461 844 462 ne
rect 844 461 909 462
tri 909 461 910 462 sw
tri 1299 461 1300 462 ne
rect 1300 461 1365 462
tri 1365 461 1366 462 sw
tri 1480 461 1481 462 ne
rect 1481 461 1609 462
tri 844 460 845 461 ne
rect 845 460 910 461
tri 910 460 911 461 sw
tri 1300 460 1301 461 ne
rect 1301 460 1366 461
tri 1366 460 1367 461 sw
tri 1481 460 1482 461 ne
rect 1482 460 1609 461
tri 845 459 846 460 ne
rect 846 459 911 460
tri 911 459 912 460 sw
tri 1301 459 1302 460 ne
rect 1302 459 1367 460
tri 1367 459 1368 460 sw
tri 1482 459 1483 460 ne
rect 1483 459 1609 460
tri 846 458 847 459 ne
rect 847 458 912 459
tri 912 458 913 459 sw
tri 1302 458 1303 459 ne
rect 1303 458 1368 459
tri 1368 458 1369 459 sw
tri 1483 458 1484 459 ne
rect 1484 458 1609 459
tri 847 457 848 458 ne
rect 848 457 913 458
tri 913 457 914 458 sw
tri 1303 457 1304 458 ne
rect 1304 457 1369 458
tri 1369 457 1370 458 sw
tri 1484 457 1485 458 ne
rect 1485 457 1609 458
tri 848 456 849 457 ne
rect 849 456 914 457
tri 914 456 915 457 sw
tri 1304 456 1305 457 ne
rect 1305 456 1370 457
tri 1370 456 1371 457 sw
tri 1485 456 1486 457 ne
rect 1486 456 1609 457
tri 849 455 850 456 ne
rect 850 455 915 456
tri 915 455 916 456 sw
tri 1305 455 1306 456 ne
rect 1306 455 1371 456
tri 1371 455 1372 456 sw
tri 1486 455 1487 456 ne
rect 1487 455 1609 456
tri 850 454 851 455 ne
rect 851 454 916 455
tri 916 454 917 455 sw
tri 1306 454 1307 455 ne
rect 1307 454 1372 455
tri 1372 454 1373 455 sw
tri 1487 454 1488 455 ne
rect 1488 454 1609 455
tri 851 453 852 454 ne
rect 852 453 917 454
tri 917 453 918 454 sw
tri 1307 453 1308 454 ne
rect 1308 453 1373 454
tri 1373 453 1374 454 sw
tri 1488 453 1489 454 ne
rect 1489 453 1609 454
tri 852 452 853 453 ne
rect 853 452 918 453
tri 918 452 919 453 sw
tri 1308 452 1309 453 ne
rect 1309 452 1374 453
tri 1374 452 1375 453 sw
tri 1489 452 1490 453 ne
rect 1490 452 1609 453
tri 853 451 854 452 ne
rect 854 451 919 452
tri 919 451 920 452 sw
tri 1309 451 1310 452 ne
rect 1310 451 1375 452
tri 1375 451 1376 452 sw
tri 1490 451 1491 452 ne
rect 1491 451 1609 452
tri 854 450 855 451 ne
rect 855 450 920 451
tri 920 450 921 451 sw
tri 1310 450 1311 451 ne
rect 1311 450 1376 451
tri 1376 450 1377 451 sw
tri 1491 450 1492 451 ne
rect 1492 450 1609 451
tri 855 449 856 450 ne
rect 856 449 921 450
tri 921 449 922 450 sw
tri 1311 449 1312 450 ne
rect 1312 449 1377 450
tri 1377 449 1378 450 sw
tri 1492 449 1493 450 ne
rect 1493 449 1609 450
tri 856 448 857 449 ne
rect 857 448 922 449
tri 922 448 923 449 sw
tri 1312 448 1313 449 ne
rect 1313 448 1378 449
tri 1378 448 1379 449 sw
tri 1493 448 1494 449 ne
rect 1494 448 1609 449
tri 857 447 858 448 ne
rect 858 447 923 448
tri 923 447 924 448 sw
tri 1313 447 1314 448 ne
rect 1314 447 1379 448
tri 1379 447 1380 448 sw
tri 1494 447 1495 448 ne
rect 1495 447 1609 448
rect 244 445 663 447
tri 858 446 859 447 ne
rect 859 446 924 447
tri 924 446 925 447 sw
tri 1314 446 1315 447 ne
rect 1315 446 1380 447
tri 1380 446 1381 447 sw
tri 1495 446 1496 447 ne
rect 1496 446 1609 447
tri 859 445 860 446 ne
rect 860 445 925 446
tri 925 445 926 446 sw
tri 1315 445 1316 446 ne
rect 1316 445 1381 446
tri 1381 445 1382 446 sw
tri 1496 445 1497 446 ne
rect 1497 445 1609 446
tri 461 430 476 445 ne
rect 476 430 663 445
tri 860 444 861 445 ne
rect 861 444 926 445
tri 926 444 927 445 sw
tri 1316 444 1317 445 ne
rect 1317 444 1382 445
tri 1382 444 1383 445 sw
tri 1497 444 1498 445 ne
rect 1498 444 1609 445
tri 861 443 862 444 ne
rect 862 443 927 444
tri 927 443 928 444 sw
tri 1317 443 1318 444 ne
rect 1318 443 1383 444
tri 1383 443 1384 444 sw
tri 1498 443 1499 444 ne
rect 1499 443 1609 444
tri 862 442 863 443 ne
rect 863 442 928 443
tri 928 442 929 443 sw
tri 1318 442 1319 443 ne
rect 1319 442 1384 443
tri 1384 442 1385 443 sw
tri 1499 442 1500 443 ne
rect 1500 442 1609 443
tri 863 441 864 442 ne
rect 864 441 929 442
tri 929 441 930 442 sw
tri 1319 441 1320 442 ne
rect 1320 441 1385 442
tri 1385 441 1386 442 sw
tri 1500 441 1501 442 ne
rect 1501 441 1609 442
tri 864 440 865 441 ne
rect 865 440 930 441
tri 930 440 931 441 sw
tri 1320 440 1321 441 ne
rect 1321 440 1386 441
tri 1386 440 1387 441 sw
tri 1501 440 1502 441 ne
rect 1502 440 1609 441
tri 865 439 866 440 ne
rect 866 439 931 440
tri 931 439 932 440 sw
tri 1321 439 1322 440 ne
rect 1322 439 1387 440
tri 1387 439 1388 440 sw
tri 1502 439 1503 440 ne
rect 1503 439 1609 440
tri 866 438 867 439 ne
rect 867 438 932 439
tri 932 438 933 439 sw
tri 1322 438 1323 439 ne
rect 1323 438 1388 439
tri 1388 438 1389 439 sw
tri 1503 438 1504 439 ne
rect 1504 438 1609 439
tri 867 437 868 438 ne
rect 868 437 933 438
tri 933 437 934 438 sw
tri 1323 437 1324 438 ne
rect 1324 437 1389 438
tri 1389 437 1390 438 sw
tri 1504 437 1505 438 ne
rect 1505 437 1609 438
tri 868 436 869 437 ne
rect 869 436 934 437
tri 934 436 935 437 sw
tri 1324 436 1325 437 ne
rect 1325 436 1390 437
tri 1390 436 1391 437 sw
tri 1505 436 1506 437 ne
rect 1506 436 1609 437
tri 869 435 870 436 ne
rect 870 435 935 436
tri 935 435 936 436 sw
tri 1325 435 1326 436 ne
rect 1326 435 1391 436
tri 1391 435 1392 436 sw
tri 1506 435 1507 436 ne
rect 1507 435 1609 436
tri 870 434 871 435 ne
rect 871 434 936 435
tri 936 434 937 435 sw
tri 1326 434 1327 435 ne
rect 1327 434 1392 435
tri 1392 434 1393 435 sw
tri 1569 434 1570 435 ne
rect 1570 434 1609 435
tri 871 433 872 434 ne
rect 872 433 937 434
tri 937 433 938 434 sw
tri 1327 433 1328 434 ne
rect 1328 433 1393 434
tri 1393 433 1394 434 sw
tri 1570 433 1571 434 ne
rect 1571 433 1609 434
tri 872 432 873 433 ne
rect 873 432 938 433
tri 938 432 939 433 sw
tri 1328 432 1329 433 ne
rect 1329 432 1394 433
tri 1394 432 1395 433 sw
tri 1571 432 1572 433 ne
rect 1572 432 1609 433
tri 873 431 874 432 ne
rect 874 431 939 432
tri 939 431 940 432 sw
tri 1329 431 1330 432 ne
rect 1330 431 1395 432
tri 1395 431 1396 432 sw
tri 1572 431 1573 432 ne
rect 1573 431 1609 432
tri 874 430 875 431 ne
rect 875 430 940 431
tri 940 430 941 431 sw
tri 1330 430 1331 431 ne
rect 1331 430 1396 431
tri 1396 430 1397 431 sw
tri 1573 430 1574 431 ne
rect 1574 430 1609 431
rect 1643 430 1649 464
rect 1909 470 1955 482
tri 476 424 482 430 ne
rect 482 424 623 430
tri 482 403 503 424 ne
rect 503 403 623 424
tri 583 396 590 403 ne
rect 590 396 623 403
rect 657 396 663 430
tri 875 429 876 430 ne
rect 876 429 941 430
tri 941 429 942 430 sw
tri 1331 429 1332 430 ne
rect 1332 429 1397 430
tri 1397 429 1398 430 sw
tri 1574 429 1575 430 ne
rect 1575 429 1649 430
tri 876 428 877 429 ne
rect 877 428 942 429
tri 942 428 943 429 sw
tri 1332 428 1333 429 ne
rect 1333 428 1398 429
tri 1398 428 1399 429 sw
tri 1575 428 1576 429 ne
rect 1576 428 1649 429
tri 877 427 878 428 ne
rect 878 427 943 428
tri 943 427 944 428 sw
tri 1333 427 1334 428 ne
rect 1334 427 1399 428
tri 1399 427 1400 428 sw
tri 1576 427 1577 428 ne
rect 1577 427 1649 428
tri 878 426 879 427 ne
rect 879 426 944 427
tri 944 426 945 427 sw
tri 1334 426 1335 427 ne
rect 1335 426 1400 427
tri 1400 426 1401 427 sw
tri 1577 426 1578 427 ne
rect 1578 426 1649 427
tri 879 425 880 426 ne
rect 880 425 945 426
tri 945 425 946 426 sw
tri 1335 425 1336 426 ne
rect 1336 425 1401 426
tri 1401 425 1402 426 sw
tri 1578 425 1579 426 ne
rect 1579 425 1649 426
tri 880 424 881 425 ne
rect 881 424 946 425
tri 946 424 947 425 sw
tri 1336 424 1337 425 ne
rect 1337 424 1402 425
tri 1402 424 1403 425 sw
tri 1579 424 1580 425 ne
rect 1580 424 1649 425
tri 881 423 882 424 ne
rect 882 423 947 424
tri 947 423 948 424 sw
tri 1337 423 1338 424 ne
rect 1338 423 1403 424
tri 1403 423 1404 424 sw
tri 1580 423 1581 424 ne
rect 1581 423 1649 424
tri 882 422 883 423 ne
rect 883 422 948 423
tri 948 422 949 423 sw
tri 1338 422 1339 423 ne
rect 1339 422 1404 423
tri 1404 422 1405 423 sw
tri 1581 422 1582 423 ne
rect 1582 422 1649 423
tri 883 421 884 422 ne
rect 884 421 949 422
tri 949 421 950 422 sw
tri 1339 421 1340 422 ne
rect 1340 421 1405 422
tri 1405 421 1406 422 sw
tri 1582 421 1583 422 ne
rect 1583 421 1649 422
tri 884 420 885 421 ne
rect 885 420 950 421
tri 950 420 951 421 sw
tri 1340 420 1341 421 ne
rect 1341 420 1406 421
tri 1406 420 1407 421 sw
tri 1583 420 1584 421 ne
rect 1584 420 1649 421
tri 885 419 886 420 ne
rect 886 419 951 420
tri 951 419 952 420 sw
tri 1341 419 1342 420 ne
rect 1342 419 1407 420
tri 1407 419 1408 420 sw
tri 1584 419 1585 420 ne
rect 1585 419 1649 420
tri 886 418 887 419 ne
rect 887 418 952 419
tri 952 418 953 419 sw
tri 1342 418 1343 419 ne
rect 1343 418 1408 419
tri 1408 418 1409 419 sw
tri 1585 418 1586 419 ne
rect 1586 418 1649 419
tri 887 417 888 418 ne
rect 888 417 953 418
tri 953 417 954 418 sw
tri 1343 417 1344 418 ne
rect 1344 417 1409 418
tri 1409 417 1410 418 sw
tri 1586 417 1587 418 ne
rect 1587 417 1649 418
tri 888 416 889 417 ne
rect 889 416 954 417
tri 954 416 955 417 sw
tri 1344 416 1345 417 ne
rect 1345 416 1410 417
tri 1410 416 1411 417 sw
tri 1587 416 1588 417 ne
rect 1588 416 1649 417
tri 889 415 890 416 ne
rect 890 415 955 416
tri 955 415 956 416 sw
tri 1345 415 1346 416 ne
rect 1346 415 1411 416
tri 1411 415 1412 416 sw
tri 1588 415 1589 416 ne
rect 1589 415 1649 416
tri 890 414 891 415 ne
rect 891 414 956 415
tri 956 414 957 415 sw
tri 1346 414 1347 415 ne
rect 1347 414 1412 415
tri 1412 414 1413 415 sw
tri 1589 414 1590 415 ne
rect 1590 414 1649 415
tri 891 413 892 414 ne
rect 892 413 957 414
tri 957 413 958 414 sw
tri 1347 413 1348 414 ne
rect 1348 413 1413 414
tri 1413 413 1414 414 sw
tri 1590 413 1591 414 ne
rect 1591 413 1649 414
tri 892 412 893 413 ne
rect 893 412 958 413
tri 958 412 959 413 sw
tri 1348 412 1349 413 ne
rect 1349 412 1414 413
tri 1414 412 1415 413 sw
tri 1591 412 1592 413 ne
rect 1592 412 1649 413
tri 893 411 894 412 ne
rect 894 411 959 412
tri 959 411 960 412 sw
tri 1349 411 1350 412 ne
rect 1350 411 1415 412
tri 1415 411 1416 412 sw
tri 1592 411 1593 412 ne
rect 1593 411 1649 412
tri 894 410 895 411 ne
rect 895 410 960 411
tri 960 410 961 411 sw
tri 1350 410 1351 411 ne
rect 1351 410 1416 411
tri 1416 410 1417 411 sw
tri 1593 410 1594 411 ne
rect 1594 410 1649 411
tri 895 409 896 410 ne
rect 896 409 961 410
tri 961 409 962 410 sw
tri 1351 409 1352 410 ne
rect 1352 409 1417 410
tri 1417 409 1418 410 sw
tri 1594 409 1595 410 ne
rect 1595 409 1649 410
tri 896 408 897 409 ne
rect 897 408 962 409
tri 962 408 963 409 sw
tri 1352 408 1353 409 ne
rect 1353 408 1418 409
tri 1418 408 1419 409 sw
tri 1595 408 1596 409 ne
rect 1596 408 1649 409
tri 897 407 898 408 ne
rect 898 407 963 408
tri 963 407 964 408 sw
tri 1353 407 1354 408 ne
rect 1354 407 1419 408
tri 1419 407 1420 408 sw
tri 1596 407 1597 408 ne
rect 1597 407 1649 408
tri 898 406 899 407 ne
rect 899 406 964 407
tri 964 406 965 407 sw
tri 1354 406 1355 407 ne
rect 1355 406 1420 407
tri 1420 406 1421 407 sw
tri 1597 406 1598 407 ne
rect 1598 406 1649 407
tri 899 405 900 406 ne
rect 900 405 965 406
tri 965 405 966 406 sw
tri 1355 405 1356 406 ne
rect 1356 405 1421 406
tri 1421 405 1422 406 sw
tri 1598 405 1599 406 ne
rect 1599 405 1649 406
tri 900 404 901 405 ne
rect 901 404 966 405
tri 966 404 967 405 sw
tri 1356 404 1357 405 ne
rect 1357 404 1422 405
tri 1422 404 1423 405 sw
tri 1599 404 1600 405 ne
rect 1600 404 1649 405
tri 901 403 902 404 ne
rect 902 403 967 404
tri 967 403 968 404 sw
tri 1357 403 1358 404 ne
rect 1358 403 1423 404
tri 1423 403 1424 404 sw
tri 1600 403 1601 404 ne
rect 1601 403 1649 404
tri 902 402 903 403 ne
rect 903 402 968 403
tri 968 402 969 403 sw
tri 1358 402 1359 403 ne
rect 1359 402 1424 403
tri 1424 402 1425 403 sw
tri 1601 402 1602 403 ne
rect 1602 402 1649 403
tri 903 401 904 402 ne
rect 904 401 969 402
tri 969 401 970 402 sw
tri 1359 401 1360 402 ne
rect 1360 401 1425 402
tri 1425 401 1426 402 sw
tri 1602 401 1603 402 ne
tri 904 400 905 401 ne
rect 905 400 970 401
tri 970 400 971 401 sw
tri 1360 400 1361 401 ne
rect 1361 400 1426 401
tri 1426 400 1427 401 sw
tri 905 399 906 400 ne
rect 906 399 971 400
tri 971 399 972 400 sw
tri 1361 399 1362 400 ne
rect 1362 399 1427 400
tri 1427 399 1428 400 sw
tri 906 398 907 399 ne
rect 907 398 972 399
tri 972 398 973 399 sw
tri 1362 398 1363 399 ne
rect 1363 398 1428 399
tri 1428 398 1429 399 sw
tri 907 397 908 398 ne
rect 908 397 973 398
tri 973 397 974 398 sw
tri 1363 397 1364 398 ne
rect 1364 397 1429 398
tri 1429 397 1430 398 sw
tri 908 396 909 397 ne
rect 909 396 974 397
tri 974 396 975 397 sw
tri 1364 396 1365 397 ne
rect 1365 396 1430 397
tri 1430 396 1431 397 sw
rect 81 390 216 396
rect 81 356 93 390
rect 127 356 165 390
rect 199 356 216 390
rect 81 350 216 356
rect 319 390 458 396
tri 590 392 594 396 ne
rect 594 392 663 396
tri 594 390 596 392 ne
rect 596 390 663 392
rect 319 356 331 390
rect 365 356 403 390
rect 437 356 458 390
tri 596 369 617 390 ne
rect 319 350 458 356
rect 617 358 663 390
rect 617 324 623 358
rect 657 324 663 358
rect 719 390 854 396
tri 909 395 910 396 ne
rect 910 395 1091 396
tri 910 394 911 395 ne
rect 911 394 1091 395
tri 911 393 912 394 ne
rect 912 393 1091 394
tri 912 392 913 393 ne
rect 913 392 1091 393
tri 1365 392 1369 396 ne
rect 1369 392 1554 396
tri 913 391 914 392 ne
rect 914 391 1091 392
tri 914 390 915 391 ne
rect 915 390 1091 391
tri 1369 390 1371 392 ne
rect 1371 390 1554 392
rect 719 356 731 390
rect 765 356 803 390
rect 837 356 854 390
tri 915 389 916 390 ne
rect 916 389 968 390
tri 916 388 917 389 ne
rect 917 388 968 389
tri 917 387 918 388 ne
rect 918 387 968 388
tri 918 386 919 387 ne
rect 919 386 968 387
tri 919 385 920 386 ne
rect 920 385 968 386
tri 920 384 921 385 ne
rect 921 384 968 385
tri 921 383 922 384 ne
rect 922 383 968 384
tri 922 382 923 383 ne
rect 923 382 968 383
tri 923 381 924 382 ne
rect 924 381 968 382
tri 924 380 925 381 ne
rect 925 380 968 381
tri 925 379 926 380 ne
rect 926 379 968 380
tri 926 378 927 379 ne
rect 927 378 968 379
tri 927 377 928 378 ne
rect 928 377 968 378
tri 928 376 929 377 ne
rect 929 376 968 377
tri 929 375 930 376 ne
rect 930 375 968 376
tri 930 374 931 375 ne
rect 931 374 968 375
tri 931 373 932 374 ne
rect 932 373 968 374
tri 932 372 933 373 ne
rect 933 372 968 373
tri 933 371 934 372 ne
rect 934 371 968 372
tri 934 370 935 371 ne
rect 935 370 968 371
tri 935 369 936 370 ne
rect 936 369 968 370
tri 936 368 937 369 ne
rect 937 368 968 369
tri 937 367 938 368 ne
rect 938 367 968 368
tri 938 366 939 367 ne
rect 939 366 968 367
tri 939 365 940 366 ne
rect 940 365 968 366
tri 940 364 941 365 ne
rect 941 364 968 365
tri 941 363 942 364 ne
rect 942 363 968 364
tri 942 362 943 363 ne
rect 943 362 968 363
tri 943 361 944 362 ne
rect 944 361 968 362
tri 944 360 945 361 ne
rect 945 360 968 361
tri 945 359 946 360 ne
rect 946 359 968 360
tri 946 358 947 359 ne
rect 947 358 968 359
tri 947 357 948 358 ne
rect 948 357 968 358
tri 948 356 949 357 ne
rect 949 356 968 357
rect 1002 356 1040 390
rect 1074 356 1091 390
tri 1371 356 1405 390 ne
rect 1405 356 1431 390
rect 1465 356 1503 390
rect 1537 356 1554 390
rect 719 350 854 356
tri 949 355 950 356 ne
rect 950 355 1091 356
tri 950 354 951 355 ne
rect 951 354 1091 355
tri 951 353 952 354 ne
rect 952 353 1091 354
tri 952 352 953 353 ne
rect 953 352 1091 353
tri 953 351 954 352 ne
rect 954 351 1091 352
tri 954 350 955 351 ne
rect 955 350 1091 351
tri 1405 350 1411 356 ne
rect 1411 350 1554 356
rect 1603 392 1649 402
rect 1603 358 1609 392
rect 1643 358 1649 392
rect 1603 346 1649 358
rect 1696 435 1742 452
rect 1696 401 1702 435
rect 1736 401 1742 435
rect 1696 363 1742 401
rect 617 312 663 324
rect 1696 329 1702 363
rect 1736 329 1742 363
rect 1909 436 1915 470
rect 1949 436 1955 470
rect 1909 398 1955 436
rect 1909 364 1915 398
rect 1949 364 1955 398
rect 1909 352 1955 364
rect 1996 470 2042 482
rect 2743 478 3081 484
rect 1996 436 2002 470
rect 2036 436 2042 470
tri 3035 463 3050 478 ne
rect 3050 463 3081 478
rect 3115 463 3121 497
tri 3050 447 3066 463 ne
rect 3066 447 3121 463
rect 1996 398 2042 436
rect 1996 364 2002 398
rect 2036 364 2042 398
rect 1996 352 2042 364
rect 2173 435 2219 447
rect 2173 401 2179 435
rect 2213 401 2219 435
rect 2173 363 2219 401
tri 1742 329 1760 347 sw
tri 2155 329 2173 347 se
rect 2173 329 2179 363
rect 2213 329 2219 363
rect 1696 317 1760 329
tri 1760 317 1772 329 sw
tri 2143 317 2155 329 se
rect 2155 317 2219 329
rect 2439 435 2485 447
rect 2610 442 2662 447
rect 2439 401 2445 435
rect 2479 401 2485 435
rect 2439 363 2485 401
rect 2439 329 2445 363
rect 2479 329 2485 363
rect 2439 317 2485 329
rect 2613 435 2659 442
rect 2613 401 2619 435
rect 2653 401 2659 435
rect 2613 363 2659 401
rect 2613 329 2619 363
rect 2653 329 2659 363
rect 2613 321 2659 329
rect 2893 435 2939 447
tri 3066 444 3069 447 ne
rect 3069 437 3121 447
rect 2893 401 2899 435
rect 2933 401 2939 435
rect 2893 363 2939 401
rect 3075 425 3121 437
rect 3075 391 3081 425
rect 3115 391 3121 425
rect 3075 379 3121 391
rect 2893 329 2899 363
rect 2933 329 2939 363
rect 2610 317 2662 321
rect 2893 317 2939 329
rect 1696 313 1772 317
tri 1772 313 1776 317 sw
tri 2139 313 2143 317 se
rect 2143 313 2219 317
rect 1696 267 2219 313
rect 41 82 2632 239
rect 41 70 3225 82
rect 41 36 83 70
rect 117 36 155 70
rect 189 36 227 70
rect 261 36 299 70
rect 333 36 371 70
rect 405 36 443 70
rect 477 36 515 70
rect 549 36 587 70
rect 621 36 659 70
rect 693 36 731 70
rect 765 36 803 70
rect 837 36 875 70
rect 909 36 947 70
rect 981 36 1019 70
rect 1053 36 1091 70
rect 1125 36 1163 70
rect 1197 36 1235 70
rect 1269 36 1307 70
rect 1341 36 1379 70
rect 1413 36 1451 70
rect 1485 36 1523 70
rect 1557 36 1595 70
rect 1629 36 1667 70
rect 1701 36 1739 70
rect 1773 36 1811 70
rect 1845 36 1883 70
rect 1917 36 1955 70
rect 1989 36 2027 70
rect 2061 36 2099 70
rect 2133 36 2171 70
rect 2205 36 2243 70
rect 2277 36 2315 70
rect 2349 36 2387 70
rect 2421 36 2459 70
rect 2493 36 2531 70
rect 2565 36 2603 70
rect 2637 36 2675 70
rect 2709 36 2747 70
rect 2781 36 2819 70
rect 2853 36 2891 70
rect 2925 36 2963 70
rect 2997 36 3035 70
rect 3069 36 3107 70
rect 3141 36 3179 70
rect 3213 36 3225 70
rect 41 24 3225 36
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1663361622
transform 1 0 1452 0 1 0
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1663361622
transform -1 0 820 0 1 0
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1663361622
transform 1 0 2922 0 1 0
box -46 24 399 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1663361622
transform -1 0 2287 0 1 0
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1663361622
transform 1 0 2105 0 1 0
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1663361622
transform -1 0 1634 0 1 0
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1663361622
transform 1 0 638 0 1 0
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2v2  sky130_fd_io__hvsbt_nand2v2_0
timestamp 1663361622
transform 1 0 0 0 1 0
box -34 24 569 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1663361622
transform -1 0 3104 0 1 0
box 0 24 534 1116
<< labels >>
flabel metal1 s 1709 373 1728 393 0 FreeSans 280 90 0 0 INP_DIS_I_H_N
port 1 nsew
flabel metal1 s 1619 395 1633 412 0 FreeSans 280 90 0 0 INP_DIS_I_H
port 2 nsew
flabel metal1 s 1256 629 1302 764 0 FreeSans 280 90 0 0 INP_DIS_H_N
port 3 nsew
flabel metal1 s 719 350 854 396 0 FreeSans 280 0 0 0 DM_H_N[2]
port 4 nsew
flabel metal1 s 81 350 216 396 0 FreeSans 280 0 0 0 DM_H_N[1]
port 5 nsew
flabel metal1 s 394 380 394 380 0 FreeSans 280 0 0 0 DM_H_N[0]
port 6 nsew
flabel metal1 s 2450 414 2472 439 3 FreeSans 520 90 0 0 IB_MODE_SEL_H_N
port 7 nsew
flabel metal1 s 726 896 942 1017 3 FreeSans 520 0 0 0 VDDIO_Q
port 8 nsew
flabel metal1 s 589 65 759 172 3 FreeSans 520 0 0 0 VSSD
port 9 nsew
flabel metal1 s 2908 383 2925 408 3 FreeSans 520 90 0 0 VTRIP_SEL_H_N
port 10 nsew
flabel metal1 s 2618 345 2650 385 3 FreeSans 520 90 0 0 MODE_NORMAL_N
port 11 nsew
flabel metal1 s 2013 418 2029 472 3 FreeSans 520 90 0 0 MODE_VCCHIB_N
port 12 nsew
flabel metal1 s 3085 446 3110 499 3 FreeSans 520 90 0 0 TRIPSEL_I_H
port 13 nsew
flabel metal1 s 3129 796 3197 815 3 FreeSans 520 180 0 0 TRIPSEL_I_H_N
port 14 nsew
flabel metal1 s 1917 396 1944 435 3 FreeSans 520 90 0 0 IB_MODE_SEL_H
port 15 nsew
<< properties >>
string GDS_END 45115064
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 45092100
<< end >>
