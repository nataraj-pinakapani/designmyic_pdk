magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 36 54 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel  s 39 51 80 54 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel  s 0 46 52 49 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel  s 54 46 80 49 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel  s 62 -2 63 -1 8 ANALOG_EN
port 22 nsew signal input
rlabel 
 s 46 -2 46 35 6 ANALOG_POL
port 26 nsew signal input
rlabel � s 31 -2 31 0 8 ANALOG_SEL
port 23 nsew signal input
rlabel � s 28 -2 29 2 8 DM[2]
port 6 nsew signal input
rlabel � s 67 -2 67 -1 8 DM[1]
port 7 nsew signal input
rlabel � s 50 -2 50 -1 8 DM[0]
port 8 nsew signal input
rlabel � s 35 -2 36 0 8 ENABLE_H
port 13 nsew signal input
rlabel � s 38 -2 39 1 8 ENABLE_INP_H
port 15 nsew signal input
rlabel � s 13 -2 13 3 8 ENABLE_VDDA_H
port 14 nsew signal input
rlabel 
 s 79 -2 79 183 6 ENABLE_VDDIO
port 24 nsew signal input
rlabel � s 16 -2 17 0 8 ENABLE_VSWITCH_H
port 25 nsew signal input
rlabel � s 32 -2 32 1 8 HLD_H_N
port 9 nsew signal input
rlabel � s 27 -2 27 1 8 HLD_OVR
port 21 nsew signal input
rlabel � s 5 -2 6 2 8 IB_MODE_SEL
port 12 nsew signal input
rlabel 
 s 79 -2 80 188 6 IN
port 10 nsew signal output
rlabel 
 s 0 -2 1 176 4 IN_H
port 1 nsew signal output
rlabel � s 45 -2 46 3 8 INP_DIS
port 11 nsew signal input
rlabel � s 3 -2 4 2 8 OE_N
port 16 nsew signal input
rlabel � s 22 -2 23 4 6 OUT
port 27 nsew signal input
rlabel  s 11 103 74 165 6 PAD
port 5 nsew signal bidirectional
rlabel � s 76 -2 77 0 8 PAD_A_ESD_0_H
port 3 nsew signal bidirectional
rlabel � s 68 -2 69 0 8 PAD_A_ESD_1_H
port 4 nsew signal bidirectional
rlabel 
 s 63 -2 64 8 6 PAD_A_NOESD_H
port 2 nsew signal bidirectional
rlabel � s 78 -2 78 -1 8 SLOW
port 19 nsew signal input
rlabel � s 79 -2 79 -1 8 TIE_HI_ESD
port 17 nsew signal output
rlabel � s 80 -2 80 176 6 TIE_LO_ESD
port 18 nsew signal output
rlabel  s 0 7 1 11 4 VCCD
port 36 nsew power bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 36 nsew power bidirectional
rlabel  s 79 7 80 11 6 VCCD
port 36 nsew power bidirectional
rlabel  s 79 7 80 12 6 VCCD
port 36 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 34 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 34 nsew power bidirectional
rlabel  s 79 0 80 5 6 VCCHIB
port 34 nsew power bidirectional
rlabel  s 79 0 80 5 6 VCCHIB
port 34 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 31 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 31 nsew power bidirectional
rlabel  s 79 13 80 16 6 VDDA
port 31 nsew power bidirectional
rlabel  s 79 13 80 16 6 VDDA
port 31 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 68 80 93 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 18 80 22 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 18 80 22 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 68 80 93 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 79 62 80 66 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 79 62 80 67 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 46 3 46 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 54 3 55 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 46 80 55 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 35 80 38 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 50 80 51 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 47 54 80 55 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 47 46 80 46 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 35 80 38 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 38 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 38 nsew ground bidirectional
rlabel  s 79 40 80 44 6 VSSD
port 38 nsew ground bidirectional
rlabel  s 79 40 80 44 6 VSSD
port 38 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 174 80 198 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 24 80 28 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 24 80 28 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 174 80 198 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 79 56 80 61 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 79 56 80 61 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 32 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 32 nsew power bidirectional
rlabel  s 79 30 80 33 6 VSWITCH
port 32 nsew power bidirectional
rlabel  s 79 30 80 33 6 VSWITCH
port 32 nsew power bidirectional
rlabel � s 6 -2 6 0 8 VTRIP_SEL
port 20 nsew signal input
<< properties >>
string LEFclass PAD INOUT
string FIXED_BBOX 0 0 80 198
string LEFview TRUE
<< end >>
