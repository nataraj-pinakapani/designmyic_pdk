magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 5 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 5 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 46 5 55 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 54 5 55 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 46 5 46 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 35 5 38 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 35 5 38 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 13 5 16 6 VDDA
port 4 nsew power bidirectional
rlabel  s 0 13 5 16 6 VDDA
port 4 nsew power bidirectional
rlabel  s 0 30 5 33 6 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 30 5 33 6 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 62 5 66 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 62 5 67 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 0 5 5 6 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 0 5 5 6 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 68 5 93 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 68 5 93 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 18 5 22 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 18 5 22 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 7 5 11 6 VCCD
port 9 nsew power bidirectional
rlabel  s 0 7 5 12 6 VCCD
port 9 nsew power bidirectional
rlabel  s 0 24 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 5 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 40 5 44 6 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 40 5 44 6 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 56 5 61 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 56 5 61 6 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string LEFclass PAD SPACER
string FIXED_BBOX 0 0 5 198
string LEFview TRUE
<< end >>
