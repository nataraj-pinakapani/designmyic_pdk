magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -1149 1466 -818 1530
rect -1515 1427 -744 1466
rect -1515 728 -692 1427
rect -1258 727 -692 728
rect 8626 697 9486 1429
rect -1516 -706 -730 -540
<< pwell >>
rect -1407 2496 -807 2582
rect 8774 1597 9446 1849
rect -1172 566 -894 622
rect -1452 563 -894 566
rect -1618 430 -894 563
rect -1618 160 -1474 430
<< mvnmos >>
rect 8867 1623 8987 1823
rect 9043 1623 9163 1823
rect 9247 1623 9367 1823
rect -1373 456 -1273 540
rect -1093 456 -973 596
<< mvpmos >>
rect -1373 794 -1273 1394
rect -1093 1062 -973 1262
rect -1093 794 -973 994
rect 8867 763 8987 1363
rect 9043 763 9163 1363
rect 9247 763 9367 1363
<< mvndiff >>
rect 8800 1805 8867 1823
rect 8800 1771 8808 1805
rect 8842 1771 8867 1805
rect 8800 1737 8867 1771
rect 8800 1703 8808 1737
rect 8842 1703 8867 1737
rect 8800 1669 8867 1703
rect 8800 1635 8808 1669
rect 8842 1635 8867 1669
rect 8800 1623 8867 1635
rect 8987 1805 9043 1823
rect 8987 1771 8998 1805
rect 9032 1771 9043 1805
rect 8987 1737 9043 1771
rect 8987 1703 8998 1737
rect 9032 1703 9043 1737
rect 8987 1669 9043 1703
rect 8987 1635 8998 1669
rect 9032 1635 9043 1669
rect 8987 1623 9043 1635
rect 9163 1805 9247 1823
rect 9163 1771 9188 1805
rect 9222 1771 9247 1805
rect 9163 1737 9247 1771
rect 9163 1703 9188 1737
rect 9222 1703 9247 1737
rect 9163 1669 9247 1703
rect 9163 1635 9188 1669
rect 9222 1635 9247 1669
rect 9163 1623 9247 1635
rect 9367 1805 9420 1823
rect 9367 1771 9378 1805
rect 9412 1771 9420 1805
rect 9367 1737 9420 1771
rect 9367 1703 9378 1737
rect 9412 1703 9420 1737
rect 9367 1669 9420 1703
rect 9367 1635 9378 1669
rect 9412 1635 9420 1669
rect 9367 1623 9420 1635
rect -1146 584 -1093 596
rect -1146 550 -1138 584
rect -1104 550 -1093 584
rect -1426 528 -1373 540
rect -1426 494 -1418 528
rect -1384 494 -1373 528
rect -1426 456 -1373 494
rect -1273 528 -1220 540
rect -1273 494 -1262 528
rect -1228 494 -1220 528
rect -1273 456 -1220 494
rect -1146 516 -1093 550
rect -1146 482 -1138 516
rect -1104 482 -1093 516
rect -1146 456 -1093 482
rect -973 584 -920 596
rect -973 550 -962 584
rect -928 550 -920 584
rect -973 516 -920 550
rect -973 482 -962 516
rect -928 482 -920 516
rect -973 456 -920 482
<< mvpdiff >>
rect -1426 1382 -1373 1394
rect -1426 1348 -1418 1382
rect -1384 1348 -1373 1382
rect -1426 1314 -1373 1348
rect -1426 1280 -1418 1314
rect -1384 1280 -1373 1314
rect -1426 1246 -1373 1280
rect -1426 1212 -1418 1246
rect -1384 1212 -1373 1246
rect -1426 1178 -1373 1212
rect -1426 1144 -1418 1178
rect -1384 1144 -1373 1178
rect -1426 1110 -1373 1144
rect -1426 1076 -1418 1110
rect -1384 1076 -1373 1110
rect -1426 1042 -1373 1076
rect -1426 1008 -1418 1042
rect -1384 1008 -1373 1042
rect -1426 974 -1373 1008
rect -1426 940 -1418 974
rect -1384 940 -1373 974
rect -1426 906 -1373 940
rect -1426 872 -1418 906
rect -1384 872 -1373 906
rect -1426 794 -1373 872
rect -1273 1382 -1220 1394
rect -1273 1348 -1262 1382
rect -1228 1348 -1220 1382
rect -1273 1314 -1220 1348
rect -1273 1280 -1262 1314
rect -1228 1280 -1220 1314
rect -1273 1246 -1220 1280
rect -1273 1212 -1262 1246
rect -1228 1212 -1220 1246
rect -1273 1178 -1220 1212
rect -1273 1144 -1262 1178
rect -1228 1144 -1220 1178
rect -1273 1110 -1220 1144
rect -1273 1076 -1262 1110
rect -1228 1076 -1220 1110
rect -1273 1042 -1220 1076
rect -1146 1244 -1093 1262
rect -1146 1210 -1138 1244
rect -1104 1210 -1093 1244
rect -1146 1176 -1093 1210
rect -1146 1142 -1138 1176
rect -1104 1142 -1093 1176
rect -1146 1108 -1093 1142
rect -1146 1074 -1138 1108
rect -1104 1074 -1093 1108
rect -1146 1062 -1093 1074
rect -973 1244 -920 1262
rect -973 1210 -962 1244
rect -928 1210 -920 1244
rect -973 1176 -920 1210
rect -973 1142 -962 1176
rect -928 1142 -920 1176
rect -973 1108 -920 1142
rect -973 1074 -962 1108
rect -928 1074 -920 1108
rect -973 1062 -920 1074
rect -1273 1008 -1262 1042
rect -1228 1008 -1220 1042
rect -1273 974 -1220 1008
rect -1273 940 -1262 974
rect -1228 940 -1220 974
rect -1273 906 -1220 940
rect -1273 872 -1262 906
rect -1228 872 -1220 906
rect -1273 794 -1220 872
rect -1146 982 -1093 994
rect -1146 948 -1138 982
rect -1104 948 -1093 982
rect -1146 914 -1093 948
rect -1146 880 -1138 914
rect -1104 880 -1093 914
rect -1146 846 -1093 880
rect -1146 812 -1138 846
rect -1104 812 -1093 846
rect -1146 794 -1093 812
rect -973 982 -920 994
rect -973 948 -962 982
rect -928 948 -920 982
rect -973 914 -920 948
rect -973 880 -962 914
rect -928 880 -920 914
rect -973 846 -920 880
rect -973 812 -962 846
rect -928 812 -920 846
rect -973 794 -920 812
rect 8800 1351 8867 1363
rect 8800 1317 8808 1351
rect 8842 1317 8867 1351
rect 8800 1283 8867 1317
rect 8800 1249 8808 1283
rect 8842 1249 8867 1283
rect 8800 1215 8867 1249
rect 8800 1181 8808 1215
rect 8842 1181 8867 1215
rect 8800 1147 8867 1181
rect 8800 1113 8808 1147
rect 8842 1113 8867 1147
rect 8800 1079 8867 1113
rect 8800 1045 8808 1079
rect 8842 1045 8867 1079
rect 8800 1011 8867 1045
rect 8800 977 8808 1011
rect 8842 977 8867 1011
rect 8800 943 8867 977
rect 8800 909 8808 943
rect 8842 909 8867 943
rect 8800 875 8867 909
rect 8800 841 8808 875
rect 8842 841 8867 875
rect 8800 763 8867 841
rect 8987 763 9043 1363
rect 9163 1351 9247 1363
rect 9163 1317 9188 1351
rect 9222 1317 9247 1351
rect 9163 1283 9247 1317
rect 9163 1249 9188 1283
rect 9222 1249 9247 1283
rect 9163 1215 9247 1249
rect 9163 1181 9188 1215
rect 9222 1181 9247 1215
rect 9163 1147 9247 1181
rect 9163 1113 9188 1147
rect 9222 1113 9247 1147
rect 9163 1079 9247 1113
rect 9163 1045 9188 1079
rect 9222 1045 9247 1079
rect 9163 1011 9247 1045
rect 9163 977 9188 1011
rect 9222 977 9247 1011
rect 9163 943 9247 977
rect 9163 909 9188 943
rect 9222 909 9247 943
rect 9163 875 9247 909
rect 9163 841 9188 875
rect 9222 841 9247 875
rect 9163 763 9247 841
rect 9367 1351 9420 1363
rect 9367 1317 9378 1351
rect 9412 1317 9420 1351
rect 9367 1283 9420 1317
rect 9367 1249 9378 1283
rect 9412 1249 9420 1283
rect 9367 1215 9420 1249
rect 9367 1181 9378 1215
rect 9412 1181 9420 1215
rect 9367 1147 9420 1181
rect 9367 1113 9378 1147
rect 9412 1113 9420 1147
rect 9367 1079 9420 1113
rect 9367 1045 9378 1079
rect 9412 1045 9420 1079
rect 9367 1011 9420 1045
rect 9367 977 9378 1011
rect 9412 977 9420 1011
rect 9367 943 9420 977
rect 9367 909 9378 943
rect 9412 909 9420 943
rect 9367 875 9420 909
rect 9367 841 9378 875
rect 9412 841 9420 875
rect 9367 763 9420 841
<< mvndiffc >>
rect 8808 1771 8842 1805
rect 8808 1703 8842 1737
rect 8808 1635 8842 1669
rect 8998 1771 9032 1805
rect 8998 1703 9032 1737
rect 8998 1635 9032 1669
rect 9188 1771 9222 1805
rect 9188 1703 9222 1737
rect 9188 1635 9222 1669
rect 9378 1771 9412 1805
rect 9378 1703 9412 1737
rect 9378 1635 9412 1669
rect -1138 550 -1104 584
rect -1418 494 -1384 528
rect -1262 494 -1228 528
rect -1138 482 -1104 516
rect -962 550 -928 584
rect -962 482 -928 516
<< mvpdiffc >>
rect -1418 1348 -1384 1382
rect -1418 1280 -1384 1314
rect -1418 1212 -1384 1246
rect -1418 1144 -1384 1178
rect -1418 1076 -1384 1110
rect -1418 1008 -1384 1042
rect -1418 940 -1384 974
rect -1418 872 -1384 906
rect -1262 1348 -1228 1382
rect -1262 1280 -1228 1314
rect -1262 1212 -1228 1246
rect -1262 1144 -1228 1178
rect -1262 1076 -1228 1110
rect -1138 1210 -1104 1244
rect -1138 1142 -1104 1176
rect -1138 1074 -1104 1108
rect -962 1210 -928 1244
rect -962 1142 -928 1176
rect -962 1074 -928 1108
rect -1262 1008 -1228 1042
rect -1262 940 -1228 974
rect -1262 872 -1228 906
rect -1138 948 -1104 982
rect -1138 880 -1104 914
rect -1138 812 -1104 846
rect -962 948 -928 982
rect -962 880 -928 914
rect -962 812 -928 846
rect 8808 1317 8842 1351
rect 8808 1249 8842 1283
rect 8808 1181 8842 1215
rect 8808 1113 8842 1147
rect 8808 1045 8842 1079
rect 8808 977 8842 1011
rect 8808 909 8842 943
rect 8808 841 8842 875
rect 9188 1317 9222 1351
rect 9188 1249 9222 1283
rect 9188 1181 9222 1215
rect 9188 1113 9222 1147
rect 9188 1045 9222 1079
rect 9188 977 9222 1011
rect 9188 909 9222 943
rect 9188 841 9222 875
rect 9378 1317 9412 1351
rect 9378 1249 9412 1283
rect 9378 1181 9412 1215
rect 9378 1113 9412 1147
rect 9378 1045 9412 1079
rect 9378 977 9412 1011
rect 9378 909 9412 943
rect 9378 841 9412 875
<< psubdiff >>
rect -1592 513 -1522 537
rect -1592 479 -1563 513
rect -1529 479 -1522 513
rect -1592 423 -1522 479
rect -1592 389 -1563 423
rect -1529 389 -1522 423
rect -1592 333 -1522 389
rect -1592 299 -1563 333
rect -1529 299 -1522 333
rect -1592 244 -1522 299
rect -1592 210 -1563 244
rect -1529 210 -1522 244
rect -1592 186 -1522 210
<< mvpsubdiff >>
rect -1381 2522 -1357 2556
rect -1323 2522 -1279 2556
rect -1245 2522 -1201 2556
rect -1167 2522 -1123 2556
rect -1089 2522 -1045 2556
rect -1011 2522 -968 2556
rect -934 2522 -891 2556
rect -857 2522 -833 2556
rect -1522 186 -1500 537
<< mvnsubdiff >>
rect -1083 1430 -1059 1464
rect -1025 1430 -942 1464
rect -908 1430 -884 1464
rect 8692 1339 8726 1363
rect 8692 1265 8726 1305
rect 8692 1191 8726 1231
rect 8692 1117 8726 1157
rect 8692 1043 8726 1083
rect 8692 969 8726 1009
rect 8692 895 8726 935
rect 8692 821 8726 861
rect 8692 763 8726 787
rect -1450 -640 -1426 -606
rect -1392 -640 -1354 -606
rect -1320 -640 -1282 -606
rect -1248 -640 -1210 -606
rect -1176 -640 -1138 -606
rect -1104 -640 -1067 -606
rect -1033 -640 -996 -606
rect -962 -640 -925 -606
rect -891 -640 -854 -606
rect -820 -640 -796 -606
<< psubdiffcont >>
rect -1563 479 -1529 513
rect -1563 389 -1529 423
rect -1563 299 -1529 333
rect -1563 210 -1529 244
<< mvpsubdiffcont >>
rect -1357 2522 -1323 2556
rect -1279 2522 -1245 2556
rect -1201 2522 -1167 2556
rect -1123 2522 -1089 2556
rect -1045 2522 -1011 2556
rect -968 2522 -934 2556
rect -891 2522 -857 2556
<< mvnsubdiffcont >>
rect -1059 1430 -1025 1464
rect -942 1430 -908 1464
rect 8692 1305 8726 1339
rect 8692 1231 8726 1265
rect 8692 1157 8726 1191
rect 8692 1083 8726 1117
rect 8692 1009 8726 1043
rect 8692 935 8726 969
rect 8692 861 8726 895
rect 8692 787 8726 821
rect -1426 -640 -1392 -606
rect -1354 -640 -1320 -606
rect -1282 -640 -1248 -606
rect -1210 -640 -1176 -606
rect -1138 -640 -1104 -606
rect -1067 -640 -1033 -606
rect -996 -640 -962 -606
rect -925 -640 -891 -606
rect -854 -640 -820 -606
<< poly >>
rect 8867 1823 8987 1849
rect 9043 1823 9163 1849
rect 9247 1823 9367 1849
rect 8867 1513 8987 1623
rect 8867 1479 8910 1513
rect 8944 1479 8987 1513
rect 8867 1445 8987 1479
rect -1373 1394 -1273 1420
rect 8867 1411 8910 1445
rect 8944 1411 8987 1445
rect 8867 1363 8987 1411
rect 9043 1513 9163 1623
rect 9043 1479 9086 1513
rect 9120 1479 9163 1513
rect 9043 1445 9163 1479
rect 9043 1411 9086 1445
rect 9120 1411 9163 1445
rect 9043 1363 9163 1411
rect 9247 1513 9367 1623
rect 9247 1479 9263 1513
rect 9297 1479 9367 1513
rect 9247 1445 9367 1479
rect 9247 1411 9263 1445
rect 9297 1411 9367 1445
rect 9247 1363 9367 1411
rect -1093 1262 -973 1288
rect -1093 994 -973 1062
rect -1373 703 -1273 794
rect -1373 669 -1342 703
rect -1308 669 -1273 703
rect -1373 635 -1273 669
rect -1373 601 -1342 635
rect -1308 601 -1273 635
rect -1373 540 -1273 601
rect -1093 746 -973 794
rect -1093 712 -1049 746
rect -1015 712 -973 746
rect 8867 737 8987 763
rect 9043 737 9163 763
rect 9247 737 9367 763
rect -1093 678 -973 712
rect -1093 644 -1049 678
rect -1015 644 -973 678
rect -1093 596 -973 644
rect -1373 430 -1273 456
rect -1093 430 -973 456
<< polycont >>
rect 8910 1479 8944 1513
rect 8910 1411 8944 1445
rect 9086 1479 9120 1513
rect 9086 1411 9120 1445
rect 9263 1479 9297 1513
rect 9263 1411 9297 1445
rect -1342 669 -1308 703
rect -1342 601 -1308 635
rect -1049 712 -1015 746
rect -1049 644 -1015 678
<< locali >>
rect -1381 2522 -1371 2556
rect -1323 2522 -1292 2556
rect -1245 2522 -1213 2556
rect -1167 2522 -1135 2556
rect -1089 2522 -1057 2556
rect -1011 2522 -979 2556
rect -934 2522 -901 2556
rect -857 2522 -833 2556
rect -1311 2182 -1277 2220
rect -1131 2182 -1097 2220
rect -958 2182 -924 2220
rect -1049 1911 -1015 1949
rect -1401 1814 -1367 1852
rect 8808 1805 8842 1813
rect 8808 1737 8842 1741
rect 8808 1669 8842 1703
rect 8808 1619 8842 1635
rect 8998 1805 9032 1821
rect 8998 1737 9032 1771
rect 8998 1669 9032 1703
rect 8998 1585 9032 1635
rect 9188 1805 9222 1813
rect 9188 1737 9222 1741
rect 9188 1669 9222 1703
rect 9188 1619 9222 1635
rect 9378 1805 9412 1821
rect 9378 1737 9412 1771
rect 9378 1669 9412 1703
rect 8808 1551 9313 1585
rect -1083 1430 -1059 1464
rect -1025 1430 -998 1464
rect -964 1430 -942 1464
rect -892 1430 -884 1464
rect -1418 1382 -1384 1398
rect -1418 1314 -1384 1348
rect -1418 1246 -1384 1280
rect -1418 1184 -1384 1212
rect -1418 1112 -1384 1144
rect -1418 1042 -1384 1076
rect -1418 974 -1384 1008
rect -1418 906 -1384 940
rect -1592 503 -1586 537
rect -1552 513 -1514 537
rect -1529 503 -1514 513
rect -1592 479 -1563 503
rect -1529 479 -1480 503
rect -1592 459 -1480 479
rect -1418 528 -1384 872
rect -1262 1382 -1228 1398
rect -1262 1314 -1228 1327
rect 8692 1339 8726 1363
rect -1262 1246 -1228 1255
rect -1262 1178 -1228 1183
rect -1262 1110 -1228 1144
rect -1262 1042 -1228 1076
rect -1262 974 -1228 1008
rect -1262 906 -1228 940
rect -1262 856 -1228 872
rect 8692 1265 8726 1305
rect -1138 1244 -1104 1256
rect -1138 1176 -1104 1184
rect -1138 1108 -1104 1142
rect -1138 982 -1104 1074
rect -1138 914 -1104 948
rect -1138 846 -1104 880
rect -1138 796 -1104 812
rect -962 1244 -928 1262
rect -962 1176 -928 1210
rect -962 1108 -928 1142
rect -962 1012 -928 1074
rect 8692 1191 8726 1231
rect 8808 1351 8842 1551
rect 9247 1513 9313 1551
rect 9378 1523 9412 1635
rect 8894 1479 8910 1513
rect 8944 1479 8960 1513
rect 8894 1445 8960 1479
rect 8894 1441 8910 1445
rect 8944 1441 8960 1445
rect 9070 1479 9086 1513
rect 9120 1479 9136 1513
rect 9070 1445 9136 1479
rect 9070 1441 9086 1445
rect 8944 1411 8948 1441
rect 8910 1407 8948 1411
rect 9083 1411 9086 1441
rect 9120 1441 9136 1445
rect 9247 1479 9263 1513
rect 9297 1479 9313 1513
rect 9397 1489 9435 1523
rect 9247 1445 9313 1479
rect 9120 1411 9121 1441
rect 9083 1407 9121 1411
rect 9247 1411 9263 1445
rect 9297 1411 9313 1445
rect 8808 1283 8842 1317
rect 8808 1215 8842 1249
rect 9188 1351 9222 1367
rect 9188 1283 9222 1317
rect 9188 1215 9222 1249
rect 8842 1181 8853 1209
rect 8815 1175 8853 1181
rect 8692 1117 8726 1157
rect 8692 1043 8726 1083
rect -962 982 -819 1012
rect -928 978 -819 982
rect -928 948 -785 978
rect -962 940 -785 948
rect -962 914 -819 940
rect -928 906 -819 914
rect 8692 969 8726 1009
rect 8692 895 8726 935
rect -962 846 -928 880
rect -1049 746 -1015 751
rect -1342 705 -1308 719
rect -1342 635 -1308 669
rect -1065 679 -1049 746
rect -1015 679 -999 746
rect -1065 678 -999 679
rect -1065 644 -1049 678
rect -1015 644 -999 678
rect -1342 585 -1308 599
rect -1138 584 -1104 600
rect -1418 478 -1384 494
rect -1262 539 -1228 544
rect -1592 425 -1586 459
rect -1552 425 -1514 459
rect -1262 467 -1228 494
rect -1138 539 -1104 550
rect -1138 467 -1104 482
rect -962 584 -928 812
rect -962 516 -928 550
rect -241 616 -135 887
rect 8692 836 8726 861
rect 8808 1147 8842 1175
rect 8808 1079 8842 1113
rect 8808 1011 8842 1045
rect 8808 943 8842 977
rect 8808 875 8842 909
rect 8808 825 8842 841
rect 9188 1147 9222 1181
rect 9188 1079 9222 1113
rect 9188 1011 9222 1045
rect 9188 943 9222 977
rect 9188 875 9222 909
rect 9188 836 9222 841
rect 8692 764 8726 787
rect 9378 1351 9412 1489
rect 9378 1283 9412 1317
rect 9378 1215 9412 1249
rect 9378 1147 9412 1181
rect 9378 1079 9412 1113
rect 9378 1011 9412 1045
rect 9378 943 9412 977
rect 9378 875 9412 909
rect 9378 825 9412 841
rect 9188 764 9222 802
rect -207 582 -169 616
rect -241 493 -135 582
rect 9765 578 9803 612
rect -962 466 -928 482
rect -1592 423 -1480 425
rect -1592 389 -1563 423
rect -1529 389 -1480 423
rect -1592 381 -1480 389
rect -1592 347 -1586 381
rect -1552 347 -1514 381
rect -1592 333 -1480 347
rect -1592 304 -1563 333
rect -1529 304 -1480 333
rect -1592 270 -1586 304
rect -1529 299 -1514 304
rect -1552 270 -1514 299
rect -1592 244 -1480 270
rect -1592 227 -1563 244
rect -1529 227 -1480 244
rect -1592 193 -1586 227
rect -1529 210 -1514 227
rect -1552 193 -1514 210
rect -1592 186 -1480 193
rect -940 61 -902 95
rect -1315 18 -1281 56
rect 6259 52 6297 86
rect -1150 -30 -1084 -16
rect -1150 -64 -1125 -30
rect -1091 -64 -1084 -30
rect -1150 -102 -1084 -64
rect -1150 -113 -1125 -102
rect -1091 -113 -1084 -102
rect -1082 -217 -1044 -183
rect -1378 -381 -1340 -347
rect -1314 -606 -1263 -604
rect -1229 -606 -1178 -604
rect -1144 -606 -1093 -604
rect -1059 -606 -1008 -604
rect -974 -606 -923 -604
rect -1450 -640 -1426 -606
rect -1392 -640 -1354 -606
rect -1314 -638 -1282 -606
rect -1229 -638 -1210 -606
rect -1144 -638 -1138 -606
rect -1320 -640 -1282 -638
rect -1248 -640 -1210 -638
rect -1176 -640 -1138 -638
rect -1104 -638 -1093 -606
rect -1033 -638 -1008 -606
rect -1104 -640 -1067 -638
rect -1033 -640 -996 -638
rect -962 -640 -925 -606
rect -889 -638 -854 -606
rect -891 -640 -854 -638
rect -820 -640 -796 -606
<< viali >>
rect -1371 2522 -1357 2556
rect -1357 2522 -1337 2556
rect -1292 2522 -1279 2556
rect -1279 2522 -1258 2556
rect -1213 2522 -1201 2556
rect -1201 2522 -1179 2556
rect -1135 2522 -1123 2556
rect -1123 2522 -1101 2556
rect -1057 2522 -1045 2556
rect -1045 2522 -1023 2556
rect -979 2522 -968 2556
rect -968 2522 -945 2556
rect -901 2522 -891 2556
rect -891 2522 -867 2556
rect -1311 2220 -1277 2254
rect -1311 2148 -1277 2182
rect -1131 2220 -1097 2254
rect -1131 2148 -1097 2182
rect -958 2220 -924 2254
rect -958 2148 -924 2182
rect -1049 1949 -1015 1983
rect -1401 1852 -1367 1886
rect -1049 1877 -1015 1911
rect -1401 1780 -1367 1814
rect 8808 1813 8842 1847
rect 8808 1771 8842 1775
rect 8808 1741 8842 1771
rect 9188 1813 9222 1847
rect 9188 1771 9222 1775
rect 9188 1741 9222 1771
rect -998 1430 -964 1464
rect -926 1430 -908 1464
rect -908 1430 -892 1464
rect -1418 1178 -1384 1184
rect -1418 1150 -1384 1178
rect -1418 1110 -1384 1112
rect -1418 1078 -1384 1110
rect -1586 513 -1552 537
rect -1586 503 -1563 513
rect -1563 503 -1552 513
rect -1514 503 -1480 537
rect -1262 1348 -1228 1361
rect -1262 1327 -1228 1348
rect -1262 1280 -1228 1289
rect -1262 1255 -1228 1280
rect -1262 1212 -1228 1217
rect -1262 1183 -1228 1212
rect -1138 1256 -1104 1290
rect -1138 1210 -1104 1218
rect -1138 1184 -1104 1210
rect 8876 1407 8910 1441
rect 8948 1407 8982 1441
rect 9049 1407 9083 1441
rect 9363 1489 9397 1523
rect 9435 1489 9469 1523
rect 9121 1407 9155 1441
rect 8781 1181 8808 1209
rect 8808 1181 8815 1209
rect 8781 1175 8815 1181
rect 8853 1175 8887 1209
rect -819 978 -785 1012
rect -819 906 -785 940
rect -1049 751 -1015 785
rect -1342 703 -1308 705
rect -1342 671 -1308 703
rect -1049 712 -1015 713
rect -1049 679 -1015 712
rect -1342 601 -1308 633
rect -1342 599 -1308 601
rect -1262 528 -1228 539
rect -1262 505 -1228 528
rect -1586 425 -1552 459
rect -1514 425 -1480 459
rect -1262 433 -1228 467
rect -1138 516 -1104 539
rect -1138 505 -1104 516
rect -1138 433 -1104 467
rect 8692 821 8726 836
rect 8692 802 8726 821
rect 8692 730 8726 764
rect 9188 802 9222 836
rect 9188 730 9222 764
rect -241 582 -207 616
rect -169 582 -135 616
rect 9731 578 9765 612
rect 9803 578 9837 612
rect -1586 347 -1552 381
rect -1514 347 -1480 381
rect -1586 299 -1563 304
rect -1563 299 -1552 304
rect -1586 270 -1552 299
rect -1514 270 -1480 304
rect -1586 210 -1563 227
rect -1563 210 -1552 227
rect -1586 193 -1552 210
rect -1514 193 -1480 227
rect -1315 56 -1281 90
rect -974 61 -940 95
rect -902 61 -868 95
rect 6225 52 6259 86
rect 6297 52 6331 86
rect -1315 -16 -1281 18
rect -1125 -64 -1091 -30
rect -1125 -136 -1091 -102
rect -1116 -217 -1082 -183
rect -1044 -217 -1010 -183
rect -1412 -381 -1378 -347
rect -1340 -381 -1306 -347
rect -1348 -606 -1314 -604
rect -1263 -606 -1229 -604
rect -1178 -606 -1144 -604
rect -1093 -606 -1059 -604
rect -1008 -606 -974 -604
rect -923 -606 -889 -604
rect -1348 -638 -1320 -606
rect -1320 -638 -1314 -606
rect -1263 -638 -1248 -606
rect -1248 -638 -1229 -606
rect -1178 -638 -1176 -606
rect -1176 -638 -1144 -606
rect -1093 -638 -1067 -606
rect -1067 -638 -1059 -606
rect -1008 -638 -996 -606
rect -996 -638 -974 -606
rect -923 -638 -891 -606
rect -891 -638 -889 -606
<< metal1 >>
tri 7377 3657 7451 3731 se
rect 7451 3657 9696 3731
rect 0 3645 9696 3657
rect 0 3511 7361 3645
tri 7361 3511 7495 3645 nw
tri 8852 3611 8858 3617 se
rect 8858 3611 8864 3617
tri 7613 3565 7659 3611 se
rect 7659 3565 8864 3611
rect 8916 3565 8928 3617
rect 8980 3565 8986 3617
tri 7593 3545 7613 3565 se
rect 7613 3545 7659 3565
tri 7659 3545 7679 3565 nw
tri 7559 3511 7593 3545 se
tri 7527 3479 7559 3511 se
rect 7559 3479 7593 3511
tri 7593 3479 7659 3545 nw
tri 7498 3450 7527 3479 se
rect 7527 3450 7564 3479
tri 7564 3450 7593 3479 nw
tri 6891 3427 6914 3450 se
rect 6914 3427 7518 3450
rect 4524 3375 4530 3427
rect 4582 3375 4594 3427
rect 4646 3402 5939 3427
tri 5939 3402 5964 3427 sw
tri 6866 3402 6891 3427 se
rect 6891 3404 7518 3427
tri 7518 3404 7564 3450 nw
rect 6891 3402 6932 3404
tri 6932 3402 6934 3404 nw
rect 4646 3381 6911 3402
tri 6911 3381 6932 3402 nw
rect 4646 3375 4652 3381
tri 4652 3375 4658 3381 nw
tri 5919 3375 5925 3381 ne
rect 5925 3375 6886 3381
tri 5925 3356 5944 3375 ne
rect 5944 3356 6886 3375
tri 6886 3356 6911 3381 nw
rect 8720 3362 8726 3414
rect 8778 3362 8790 3414
rect 8842 3362 9548 3414
rect 9600 3362 9612 3414
rect 9664 3362 9670 3414
rect 9581 3196 9587 3248
rect 9639 3196 9651 3248
rect 9703 3196 9709 3248
tri 9625 3189 9632 3196 ne
rect 9632 3189 9709 3196
rect 3550 3137 3556 3189
rect 3608 3137 3620 3189
rect 3672 3137 4530 3189
rect 4582 3137 4594 3189
rect 4646 3137 4652 3189
tri 9632 3184 9637 3189 ne
rect 9637 3184 9709 3189
tri 9637 3165 9656 3184 ne
rect 9656 3170 9709 3184
tri 9709 3170 9723 3184 sw
rect 9656 3165 9723 3170
tri 9656 3155 9666 3165 ne
rect 9666 3155 9723 3165
tri 9723 3155 9738 3170 sw
tri 10816 3155 10831 3170 se
rect 10831 3164 11339 3170
rect 10831 3155 11287 3164
tri 7244 3137 7262 3155 se
rect 7262 3137 8726 3155
tri 7200 3093 7244 3137 se
rect 7244 3103 8726 3137
rect 8778 3103 8790 3155
rect 8842 3103 8848 3155
tri 9666 3152 9669 3155 ne
rect 9669 3152 9738 3155
tri 9738 3152 9741 3155 sw
tri 10813 3152 10816 3155 se
rect 10816 3152 11287 3155
tri 9669 3112 9709 3152 ne
rect 9709 3112 11287 3152
tri 9709 3108 9713 3112 ne
rect 9713 3108 11339 3112
tri 10765 3103 10770 3108 ne
rect 10770 3103 11339 3108
rect 7244 3093 7262 3103
tri 7262 3093 7272 3103 nw
tri 10770 3093 10780 3103 ne
rect 10780 3100 11339 3103
rect 10780 3093 11287 3100
tri 7186 3079 7200 3093 se
rect 7200 3079 7248 3093
tri 7248 3079 7262 3093 nw
tri 10780 3079 10794 3093 ne
rect 10794 3079 11287 3093
rect 6629 3027 6635 3079
rect 6687 3027 6699 3079
rect 6751 3027 7196 3079
tri 7196 3027 7248 3079 nw
tri 10794 3042 10831 3079 ne
rect 10831 3048 11287 3079
rect 10831 3042 11339 3048
rect 0 2833 11256 2999
rect 0 2797 851 2833
tri 851 2797 887 2833 nw
tri 1001 2797 1037 2833 ne
rect 1037 2797 11256 2833
tri 9550 2772 9575 2797 ne
rect 9575 2772 9627 2797
tri 9627 2772 9652 2797 nw
rect 9576 2770 9626 2771
rect 9575 2734 9627 2770
rect 9576 2733 9626 2734
rect 9575 2689 9627 2732
tri 10143 2714 10155 2726 se
tri 9627 2689 9652 2714 sw
tri 10118 2689 10143 2714 se
rect 10143 2689 10155 2714
rect 9575 2637 9759 2689
rect 9811 2637 9823 2689
rect 9875 2637 10202 2689
rect -1383 2556 -796 2562
rect -1383 2522 -1371 2556
rect -1337 2522 -1292 2556
rect -1258 2522 -1213 2556
rect -1179 2522 -1135 2556
rect -1101 2522 -1057 2556
rect -1023 2522 -979 2556
rect -945 2522 -901 2556
rect -867 2522 -796 2556
rect -1383 2516 -796 2522
rect -1222 2479 -1151 2488
rect -1279 2421 -960 2479
rect 0 2428 9600 2473
tri 9600 2428 9645 2473 sw
tri 9811 2428 9856 2473 se
rect 9856 2428 11256 2473
rect 0 2271 11256 2428
rect -1317 2254 -1271 2266
rect -1317 2220 -1311 2254
rect -1277 2220 -1271 2254
rect -1317 2182 -1271 2220
rect -1317 2148 -1311 2182
rect -1277 2148 -1271 2182
rect -1317 2017 -1271 2148
rect -1137 2254 -1091 2266
rect -1137 2220 -1131 2254
rect -1097 2220 -1091 2254
rect -1137 2182 -1091 2220
rect -1137 2148 -1131 2182
rect -1097 2148 -1091 2182
rect -964 2254 -918 2266
rect -964 2220 -958 2254
rect -924 2220 -918 2254
rect -964 2215 -918 2220
tri -918 2215 -890 2243 sw
rect -964 2182 -890 2215
tri -1091 2148 -1087 2152 sw
rect -964 2148 -958 2182
rect -924 2148 -890 2182
rect -1137 2136 -1087 2148
tri -1087 2136 -1075 2148 sw
rect -964 2147 -890 2148
tri -890 2147 -822 2215 sw
rect 9514 2177 9520 2229
rect 9572 2177 9584 2229
rect 9636 2215 9770 2229
tri 9770 2215 9784 2229 sw
rect 9636 2177 9784 2215
tri 9784 2177 9822 2215 sw
tri 9752 2149 9780 2177 ne
rect 9780 2150 9822 2177
tri 9822 2150 9849 2177 sw
rect 9780 2149 9934 2150
rect -964 2136 -822 2147
tri -822 2136 -811 2147 sw
rect -1137 2094 -1075 2136
tri -1075 2094 -1033 2136 sw
tri -891 2135 -890 2136 ne
rect -890 2135 -811 2136
tri -811 2135 -810 2136 sw
tri -890 2099 -854 2135 ne
rect -1137 2087 -893 2094
tri -1271 2017 -1228 2060 sw
rect -1137 2048 -945 2087
tri -993 2017 -962 2048 ne
rect -962 2035 -945 2048
rect -962 2023 -893 2035
rect -962 2017 -945 2023
rect -1317 1995 -1228 2017
tri -1228 1995 -1206 2017 sw
tri -962 2000 -945 2017 ne
rect -1317 1983 -1009 1995
rect -1317 1949 -1049 1983
rect -1015 1949 -1009 1983
rect -945 1965 -893 1971
tri -1080 1924 -1055 1949 ne
rect -1055 1911 -1009 1949
rect -1413 1892 -1361 1898
rect -1413 1826 -1361 1840
rect -1413 1768 -1361 1774
rect -1135 1887 -1083 1893
rect -1055 1877 -1049 1911
rect -1015 1877 -1009 1911
rect -1055 1865 -1009 1877
tri -886 1865 -854 1897 se
rect -854 1865 -810 2135
rect 5799 2095 5805 2147
rect 5857 2095 5869 2147
rect 5921 2145 6439 2147
tri 6439 2145 6441 2147 sw
rect 5921 2143 6441 2145
tri 6441 2143 6443 2145 sw
rect 5921 2136 6443 2143
tri 6443 2136 6450 2143 sw
rect 5921 2131 6450 2136
tri 6450 2131 6455 2136 sw
rect 5921 2095 6455 2131
tri 6417 2094 6418 2095 ne
rect 6418 2094 6455 2095
tri 6455 2094 6492 2131 sw
rect 7943 2097 7950 2149
rect 8002 2097 8014 2149
rect 8066 2147 8718 2149
tri 8718 2147 8720 2149 sw
tri 9450 2147 9452 2149 se
rect 9452 2147 9618 2149
rect 8066 2146 8720 2147
tri 8720 2146 8721 2147 sw
tri 9449 2146 9450 2147 se
rect 9450 2146 9618 2147
rect 8066 2097 9618 2146
rect 9670 2097 9682 2149
rect 9734 2097 9740 2149
tri 9780 2145 9784 2149 ne
rect 9784 2145 9934 2149
tri 9784 2131 9798 2145 ne
rect 9798 2131 9934 2145
tri 9798 2107 9822 2131 ne
rect 9822 2107 9934 2131
tri 9822 2098 9831 2107 ne
rect 9831 2098 9934 2107
rect 9986 2098 9998 2150
rect 10050 2098 10056 2150
rect 10904 2139 10956 2145
tri 10871 2098 10904 2131 se
tri 10870 2097 10871 2098 se
rect 10871 2097 10904 2098
tri 10867 2094 10870 2097 se
rect 10870 2094 10904 2097
tri 6418 2069 6443 2094 ne
rect 6443 2069 6492 2094
tri 6492 2069 6517 2094 sw
tri 10842 2069 10867 2094 se
rect 10867 2087 10904 2094
rect 10867 2075 10956 2087
rect 10867 2069 10904 2075
tri 6443 2017 6495 2069 ne
rect 6495 2017 8495 2069
rect 8547 2017 8559 2069
rect 8611 2023 10904 2069
rect 8611 2017 10956 2023
tri -892 1859 -886 1865 se
rect -886 1859 -810 1865
rect -141 1980 -89 1986
rect -141 1916 -89 1928
tri -904 1847 -892 1859 se
rect -892 1849 -810 1859
tri -143 1858 -141 1860 se
rect -141 1858 -89 1864
rect 0 1859 11256 1989
rect 11492 1907 11544 1913
tri 11486 1859 11492 1865 se
tri 8777 1858 8778 1859 ne
rect 8778 1858 9228 1859
rect -892 1847 -812 1849
tri -812 1847 -810 1849 nw
tri -154 1847 -143 1858 se
rect -143 1847 -104 1858
tri -104 1847 -93 1858 nw
tri 8778 1847 8789 1858 ne
rect 8789 1847 9228 1858
tri -911 1840 -904 1847 se
rect -904 1840 -825 1847
rect -1135 1834 -1083 1835
tri -1083 1834 -1077 1840 sw
tri -917 1834 -911 1840 se
rect -911 1834 -825 1840
tri -825 1834 -812 1847 nw
tri -167 1834 -154 1847 se
rect -154 1834 -117 1847
tri -117 1834 -104 1847 nw
tri 8789 1834 8802 1847 ne
rect -1135 1823 -1077 1834
rect -1083 1813 -1077 1823
tri -1077 1813 -1056 1834 sw
tri -938 1813 -917 1834 se
rect -917 1813 -846 1834
tri -846 1813 -825 1834 nw
tri -188 1813 -167 1834 se
rect -167 1813 -138 1834
tri -138 1813 -117 1834 nw
rect 8802 1813 8808 1847
rect 8842 1813 9188 1847
rect 9222 1813 9228 1847
tri 9228 1834 9253 1859 nw
tri 11461 1834 11486 1859 se
rect 11486 1855 11492 1859
rect 11486 1843 11544 1855
rect 11486 1834 11492 1843
tri 11458 1831 11461 1834 se
rect 11461 1831 11492 1834
rect -1083 1810 -1056 1813
tri -1056 1810 -1053 1813 sw
tri -941 1810 -938 1813 se
rect -938 1810 -849 1813
tri -849 1810 -846 1813 nw
tri -191 1810 -188 1813 se
rect -188 1810 -141 1813
tri -141 1810 -138 1813 nw
rect -1083 1775 -884 1810
tri -884 1775 -849 1810 nw
tri -226 1775 -191 1810 se
rect -191 1775 -176 1810
tri -176 1775 -141 1810 nw
rect 8802 1775 9228 1813
rect -1083 1771 -891 1775
rect -1135 1768 -891 1771
tri -891 1768 -884 1775 nw
tri -233 1768 -226 1775 se
rect -226 1768 -191 1775
rect -1135 1765 -894 1768
tri -894 1765 -891 1768 nw
tri -236 1765 -233 1768 se
rect -233 1765 -191 1768
tri -241 1760 -236 1765 se
rect -236 1760 -191 1765
tri -191 1760 -176 1775 nw
tri -245 1756 -241 1760 se
rect -241 1756 -195 1760
tri -195 1756 -191 1760 nw
tri -260 1741 -245 1756 se
rect -245 1741 -210 1756
tri -210 1741 -195 1756 nw
tri -277 1724 -260 1741 se
rect -260 1724 -227 1741
tri -227 1724 -210 1741 nw
rect 7497 1730 7875 1756
tri -291 1710 -277 1724 se
rect -277 1710 -241 1724
tri -241 1710 -227 1724 nw
tri -329 1672 -291 1710 se
rect -291 1672 -279 1710
tri -279 1672 -241 1710 nw
rect 1941 1672 1947 1724
rect 1999 1672 2011 1724
rect 2063 1708 3200 1724
tri 3200 1708 3216 1724 sw
rect 2063 1672 3216 1708
tri -341 1660 -329 1672 se
rect -329 1660 -291 1672
tri -291 1660 -279 1672 nw
tri 3178 1660 3190 1672 ne
rect 3190 1660 3216 1672
tri -344 1657 -341 1660 se
rect -341 1657 -294 1660
tri -294 1657 -291 1660 nw
tri 3190 1657 3193 1660 ne
rect 3193 1657 3216 1660
tri 3216 1657 3267 1708 sw
tri -351 1650 -344 1657 se
rect -344 1650 -301 1657
tri -301 1650 -294 1657 nw
tri 3193 1650 3200 1657 ne
rect 3200 1656 3267 1657
tri 3267 1656 3268 1657 sw
rect 6560 1656 6711 1708
rect 6763 1656 6775 1708
rect 6827 1656 7292 1708
rect 7549 1704 7875 1730
rect 7927 1704 7939 1756
rect 7991 1704 7997 1756
rect 8802 1741 8808 1775
rect 8842 1741 9188 1775
rect 9222 1741 9228 1775
rect 8802 1729 9228 1741
rect 9285 1779 9426 1831
rect 9428 1830 9464 1831
rect 9427 1780 9465 1830
rect 9428 1779 9464 1780
rect 9466 1779 9514 1831
rect 9566 1779 9578 1831
rect 9630 1779 9637 1831
tri 9637 1779 9689 1831 sw
rect 9753 1779 9759 1831
rect 9811 1779 9823 1831
rect 9875 1779 9881 1831
rect 10929 1788 10977 1820
rect 11223 1791 11492 1831
rect 11223 1785 11544 1791
rect 7549 1700 7599 1704
tri 7599 1700 7603 1704 nw
rect 7549 1678 7574 1700
rect 7497 1675 7574 1678
tri 7574 1675 7599 1700 nw
tri 9260 1675 9285 1700 se
rect 9285 1675 9337 1779
tri 9337 1754 9362 1779 nw
tri 9615 1754 9640 1779 ne
rect 9640 1754 9689 1779
tri 9640 1705 9689 1754 ne
tri 9689 1711 9757 1779 sw
tri 9804 1754 9829 1779 ne
rect 9829 1754 9881 1779
rect 9830 1752 9880 1753
rect 9830 1715 9880 1716
tri 9826 1711 9829 1714 se
rect 9829 1711 9881 1714
rect 9689 1705 9757 1711
tri 9757 1705 9763 1711 sw
tri 9820 1705 9826 1711 se
rect 9826 1705 9881 1711
tri 9689 1700 9694 1705 ne
rect 9694 1700 9763 1705
tri 9337 1675 9362 1700 sw
tri 9694 1675 9719 1700 ne
rect 9719 1689 9763 1700
tri 9763 1689 9779 1705 sw
tri 9804 1689 9820 1705 se
rect 9820 1689 9881 1705
rect 9719 1675 9881 1689
rect 7497 1666 7555 1675
rect 3200 1650 3268 1656
tri -387 1614 -351 1650 se
rect -351 1614 -341 1650
rect -1135 1574 -933 1614
tri -391 1610 -387 1614 se
rect -387 1610 -341 1614
tri -341 1610 -301 1650 nw
tri 3200 1610 3240 1650 ne
rect 3240 1628 3268 1650
tri 3268 1628 3296 1656 sw
rect 3240 1610 3296 1628
tri -394 1607 -391 1610 se
rect -391 1607 -344 1610
tri -344 1607 -341 1610 nw
tri 3240 1607 3243 1610 ne
rect 3243 1607 3296 1610
tri -427 1574 -394 1607 se
rect -394 1574 -391 1607
tri -441 1560 -427 1574 se
rect -427 1560 -391 1574
tri -391 1560 -344 1607 nw
tri -466 1535 -441 1560 se
rect -441 1535 -416 1560
tri -416 1535 -391 1560 nw
rect 244 1539 290 1607
tri 3243 1583 3267 1607 ne
rect 3267 1583 3296 1607
tri 3296 1583 3341 1628 sw
rect 6907 1623 7010 1628
tri 7010 1623 7015 1628 sw
rect 6907 1607 7015 1623
tri 7015 1607 7031 1623 sw
rect 7549 1656 7555 1666
tri 7555 1656 7574 1675 nw
rect 7549 1614 7552 1656
tri 7552 1653 7555 1656 nw
rect 8628 1623 8634 1675
rect 8686 1623 8698 1675
rect 8750 1623 9363 1675
rect 9365 1674 9401 1675
rect 9364 1624 9402 1674
rect 9365 1623 9401 1624
rect 9403 1623 9509 1675
tri 9719 1637 9757 1675 ne
rect 9757 1637 9881 1675
tri 9804 1623 9818 1637 ne
rect 9818 1623 9881 1637
rect 7497 1608 7552 1614
tri 9404 1608 9419 1623 ne
rect 9419 1612 9495 1623
tri 9495 1612 9506 1623 nw
tri 9818 1612 9829 1623 ne
rect 9419 1608 9481 1612
tri 9419 1607 9420 1608 ne
rect 9420 1607 9481 1608
rect 6907 1598 7031 1607
tri 7031 1598 7040 1607 sw
tri 9420 1598 9429 1607 ne
rect 9429 1598 9481 1607
tri 9481 1598 9495 1612 nw
tri 3267 1567 3283 1583 ne
rect 3283 1567 3556 1583
tri 244 1535 248 1539 ne
rect 248 1535 290 1539
rect -466 1529 -422 1535
tri -422 1529 -416 1535 nw
tri 248 1529 254 1535 ne
rect 254 1531 290 1535
tri 290 1531 326 1567 sw
tri 3283 1531 3319 1567 ne
rect 3319 1531 3556 1567
rect 3608 1531 3620 1583
rect 3672 1531 3678 1583
rect 6907 1576 7040 1598
tri 6988 1533 7031 1576 ne
rect 7031 1558 7040 1576
tri 7040 1558 7080 1598 sw
rect 9430 1596 9480 1597
rect 9430 1559 9480 1560
rect 7031 1533 7080 1558
tri 7080 1533 7105 1558 sw
tri 9404 1533 9429 1558 se
rect 9429 1533 9481 1558
tri 9481 1533 9506 1558 sw
tri 9804 1533 9829 1558 se
rect 9829 1533 9881 1623
tri 7031 1531 7033 1533 ne
rect 7033 1531 9561 1533
rect 254 1529 326 1531
tri 326 1529 328 1531 sw
tri 7033 1529 7035 1531 ne
rect 7035 1529 9561 1531
rect -466 1524 -427 1529
tri -427 1524 -422 1529 nw
tri 254 1524 259 1529 ne
rect 259 1524 328 1529
tri 328 1524 333 1529 sw
rect -1010 1520 -880 1524
rect -466 1523 -428 1524
tri -428 1523 -427 1524 nw
tri 259 1523 260 1524 ne
rect 260 1523 333 1524
tri 333 1523 334 1524 sw
rect 6810 1523 6862 1529
tri 7035 1524 7040 1529 ne
rect 7040 1524 9561 1529
tri 7040 1523 7041 1524 ne
rect 7041 1523 9561 1524
tri -1456 1489 -1425 1520 ne
rect -1425 1489 -650 1520
tri -1425 1464 -1400 1489 ne
rect -1400 1464 -650 1489
tri -1400 1430 -1366 1464 ne
rect -1366 1430 -998 1464
rect -964 1430 -926 1464
rect -892 1430 -650 1464
tri -1366 1407 -1343 1430 ne
rect -1343 1407 -650 1430
tri -1343 1401 -1337 1407 ne
rect -1337 1361 -650 1407
rect -1337 1327 -1262 1361
rect -1228 1327 -650 1361
rect -1337 1290 -650 1327
rect -1337 1289 -1138 1290
rect -1337 1255 -1262 1289
rect -1228 1256 -1138 1289
rect -1104 1256 -650 1290
rect -1228 1255 -650 1256
rect -1337 1218 -650 1255
rect -1337 1217 -1138 1218
rect -1424 1184 -1378 1196
rect -1424 1150 -1418 1184
rect -1384 1150 -1378 1184
rect -1337 1183 -1262 1217
rect -1228 1184 -1138 1217
rect -1104 1184 -650 1218
rect -1228 1183 -650 1184
rect -1337 1169 -650 1183
tri -479 1175 -466 1188 se
rect -466 1175 -430 1523
tri -430 1521 -428 1523 nw
tri 260 1521 262 1523 ne
rect 262 1521 334 1523
tri 262 1493 290 1521 ne
rect 290 1493 334 1521
tri 290 1489 294 1493 ne
rect 294 1489 334 1493
tri 334 1489 368 1523 sw
tri 294 1455 328 1489 ne
rect 328 1481 368 1489
tri 368 1481 376 1489 sw
tri 6803 1481 6810 1488 se
rect 328 1455 376 1481
tri 376 1455 402 1481 sw
tri 6777 1455 6803 1481 se
rect 6803 1471 6810 1481
tri 7041 1489 7075 1523 ne
rect 7075 1489 9363 1523
rect 9397 1489 9435 1523
rect 9469 1489 9561 1523
tri 7075 1488 7076 1489 ne
rect 7076 1488 9561 1489
tri 6862 1481 6869 1488 sw
tri 7076 1481 7083 1488 ne
rect 7083 1481 9561 1488
rect 9562 1482 9563 1532
rect 9599 1482 9600 1532
rect 9601 1481 9881 1533
rect 6862 1471 6869 1481
rect 6803 1459 6869 1471
rect 6803 1455 6810 1459
tri 328 1441 342 1455 ne
rect 342 1441 1172 1455
tri 342 1407 376 1441 ne
rect 376 1407 1172 1441
tri 376 1403 380 1407 ne
rect 380 1403 1172 1407
rect 1224 1403 1236 1455
rect 1288 1403 1294 1455
tri 6775 1453 6777 1455 se
rect 6777 1453 6810 1455
rect 6031 1401 6037 1453
rect 6089 1401 6101 1453
rect 6153 1407 6810 1453
rect 6862 1453 6869 1459
tri 6869 1453 6897 1481 sw
rect 6862 1407 7283 1453
rect 6153 1401 7283 1407
rect 7335 1401 7347 1453
rect 7399 1401 7405 1453
rect 8720 1401 8726 1453
rect 8778 1401 8790 1453
rect 8842 1441 8994 1453
rect 8842 1407 8876 1441
rect 8910 1407 8948 1441
rect 8982 1407 8994 1441
rect 8842 1401 8994 1407
rect 9034 1401 9040 1453
rect 9092 1401 9104 1453
rect 9156 1401 9167 1453
rect 272 1243 11256 1373
tri 8559 1209 8565 1215 se
rect 8565 1209 8899 1215
tri 8525 1175 8559 1209 se
rect 8559 1175 8781 1209
rect 8815 1175 8853 1209
rect 8887 1175 8899 1209
rect 10663 1190 11339 1196
tri -483 1171 -479 1175 se
rect -479 1174 -430 1175
rect -479 1171 -433 1174
tri -433 1171 -430 1174 nw
tri 8521 1171 8525 1175 se
rect 8525 1171 8899 1175
tri -485 1169 -483 1171 se
rect -483 1169 -452 1171
tri -502 1152 -485 1169 se
rect -485 1152 -452 1169
tri -452 1152 -433 1171 nw
tri 8502 1152 8521 1171 se
rect 8521 1169 8899 1171
rect 8942 1171 8994 1177
rect 8521 1152 8565 1169
tri 8565 1152 8582 1169 nw
rect -1424 1141 -1378 1150
tri -511 1143 -502 1152 se
rect -502 1143 -463 1152
tri -1378 1141 -1376 1143 sw
tri -513 1141 -511 1143 se
rect -511 1141 -463 1143
tri -463 1141 -452 1152 nw
tri 8491 1141 8502 1152 se
rect 8502 1141 8554 1152
tri 8554 1141 8565 1152 nw
tri 8936 1141 8942 1147 se
rect -1424 1138 -1376 1141
tri -1376 1138 -1373 1141 sw
tri -516 1138 -513 1141 se
rect -513 1138 -466 1141
tri -466 1138 -463 1141 nw
rect -1424 1112 -1373 1138
rect -1424 1078 -1418 1112
rect -1384 1102 -1373 1112
tri -1373 1102 -1337 1138 sw
tri -552 1102 -516 1138 se
rect -516 1102 -502 1138
tri -502 1102 -466 1138 nw
rect -1384 1089 -515 1102
tri -515 1089 -502 1102 nw
rect 1166 1089 1172 1141
rect 1224 1089 1236 1141
rect 1288 1089 6037 1141
rect 6089 1089 6101 1141
rect 6153 1089 6159 1141
tri 7920 1125 7936 1141 se
rect 7936 1125 8502 1141
rect -1384 1078 -531 1089
rect -1424 1073 -531 1078
tri -531 1073 -515 1089 nw
rect 6256 1073 6262 1125
rect 6314 1073 6326 1125
rect 6378 1096 7255 1125
tri 7255 1096 7284 1125 sw
tri 7891 1096 7920 1125 se
rect 7920 1096 8502 1125
rect 6378 1079 7284 1096
tri 7284 1079 7301 1096 sw
tri 7874 1079 7891 1096 se
rect 7891 1089 8502 1096
tri 8502 1089 8554 1141 nw
tri 8904 1109 8936 1141 se
rect 8936 1119 8942 1141
rect 10663 1150 11287 1190
rect 8936 1109 8994 1119
tri 11225 1116 11259 1150 ne
rect 11259 1138 11287 1150
rect 11259 1126 11339 1138
rect 11259 1116 11287 1126
tri 8672 1089 8692 1109 se
rect 8692 1107 8994 1109
rect 8692 1089 8942 1107
rect 7891 1079 7936 1089
tri 7936 1079 7946 1089 nw
tri 8662 1079 8672 1089 se
rect 8672 1079 8942 1089
rect 6378 1073 7301 1079
rect -1424 1066 -538 1073
tri -538 1066 -531 1073 nw
tri 7233 1066 7240 1073 ne
rect 7240 1066 7301 1073
tri 7240 1024 7282 1066 ne
rect 7282 1024 7301 1066
rect -827 1018 -775 1024
tri 7282 1022 7284 1024 ne
rect 7284 1022 7301 1024
tri 7301 1022 7358 1079 sw
tri 7817 1022 7874 1079 se
rect 7874 1022 7879 1079
tri 7879 1022 7936 1079 nw
tri 8638 1055 8662 1079 se
rect 8662 1071 8942 1079
rect 8662 1055 8692 1071
tri 8692 1055 8708 1071 nw
tri 8920 1055 8936 1071 ne
rect 8936 1055 8942 1071
rect 9671 1064 9677 1116
rect 9729 1064 9741 1116
rect 9793 1064 10052 1116
tri 11259 1088 11287 1116 ne
rect 11287 1068 11339 1074
tri 8632 1049 8638 1055 se
rect 8638 1049 8686 1055
tri 8686 1049 8692 1055 nw
tri 8936 1049 8942 1055 ne
rect 8942 1049 8994 1055
tri 8605 1022 8632 1049 se
rect 8632 1022 8646 1049
rect -1413 973 -1361 979
rect -1413 909 -1361 921
tri 7284 997 7309 1022 ne
rect 7309 997 7827 1022
tri -775 991 -769 997 sw
tri 7309 991 7315 997 ne
rect 7315 991 7827 997
rect -775 966 -769 991
rect -827 952 -769 966
rect -775 940 -769 952
tri -769 940 -718 991 sw
rect -775 910 -595 940
tri -595 910 -565 940 sw
rect -775 900 -565 910
tri -1361 894 -1355 900 sw
rect -827 894 -565 900
tri -565 894 -549 910 sw
rect -1361 875 -1355 894
tri -1355 875 -1336 894 sw
tri -615 875 -596 894 ne
rect -596 875 -549 894
tri -549 875 -530 894 sw
rect -1361 857 -1336 875
rect -1413 851 -1336 857
tri -1361 836 -1346 851 ne
rect -1346 848 -1336 851
tri -1336 848 -1309 875 sw
tri -596 856 -577 875 ne
rect -577 856 -530 875
tri -530 856 -511 875 sw
rect -1061 848 -624 856
tri -624 848 -616 856 sw
tri -577 848 -569 856 ne
rect -569 848 -511 856
tri -511 848 -503 856 sw
rect -1346 836 -1309 848
tri -1309 836 -1297 848 sw
rect -1061 847 -616 848
tri -616 847 -615 848 sw
tri -569 847 -568 848 ne
rect -568 847 -503 848
rect -1061 844 -615 847
tri -615 844 -612 847 sw
tri -568 844 -565 847 ne
rect -565 844 -503 847
tri -503 844 -499 848 sw
rect -1061 836 -612 844
tri -612 836 -604 844 sw
tri -565 836 -557 844 ne
rect -557 836 -499 844
tri -499 836 -491 844 sw
tri -1346 826 -1336 836 ne
rect -1336 826 -1297 836
tri -1297 826 -1287 836 sw
rect -1061 828 -604 836
tri -604 828 -596 836 sw
tri -557 828 -549 836 ne
rect -549 828 -491 836
tri -491 828 -483 836 sw
rect -1061 826 -596 828
tri -596 826 -594 828 sw
tri -549 826 -547 828 ne
rect -547 826 -483 828
tri -483 826 -481 828 sw
tri -1336 802 -1312 826 ne
rect -1312 802 -1287 826
tri -1287 802 -1263 826 sw
rect -1061 810 -594 826
rect -1061 802 -978 810
tri -978 802 -970 810 nw
tri -644 802 -636 810 ne
rect -636 802 -594 810
tri -594 802 -570 826 sw
tri -547 802 -523 826 ne
rect -523 805 -481 826
tri -481 805 -460 826 sw
rect -523 802 -460 805
tri -460 802 -457 805 sw
tri -293 802 -290 805 se
rect -290 802 -244 991
tri -1312 785 -1295 802 ne
rect -1295 785 -1263 802
tri -1263 785 -1246 802 sw
rect -1061 797 -983 802
tri -983 797 -978 802 nw
tri -636 797 -631 802 ne
rect -631 797 -570 802
tri -570 797 -565 802 sw
tri -523 797 -518 802 ne
rect -518 797 -457 802
tri -457 797 -452 802 sw
tri -298 797 -293 802 se
rect -293 797 -244 802
rect -1061 795 -999 797
tri -1295 777 -1287 785 ne
rect -1287 777 -1246 785
tri -1246 777 -1238 785 sw
tri -1287 766 -1276 777 ne
rect -1276 766 -1238 777
tri -1276 762 -1272 766 ne
rect -1411 711 -1302 717
rect -1359 705 -1302 711
rect -1359 671 -1342 705
rect -1308 671 -1302 705
rect -1359 659 -1302 671
rect -1411 645 -1302 659
rect -1359 633 -1302 645
rect -1359 599 -1342 633
rect -1308 599 -1302 633
rect -1272 679 -1238 766
rect -1061 743 -1051 795
tri -999 781 -983 797 nw
tri -631 781 -615 797 ne
rect -615 781 -565 797
tri -615 780 -614 781 ne
rect -614 780 -565 781
rect -1061 731 -999 743
tri -1238 679 -1234 683 sw
rect -1061 679 -1051 731
rect -1272 669 -1234 679
tri -1234 669 -1224 679 sw
tri -1272 621 -1224 669 ne
tri -1224 667 -1222 669 sw
rect -1061 667 -999 679
rect -809 774 -757 780
tri -614 771 -605 780 ne
rect -605 778 -565 780
tri -565 778 -546 797 sw
tri -518 778 -499 797 ne
rect -499 778 -452 797
tri -452 778 -433 797 sw
tri -317 778 -298 797 se
rect -298 779 -244 797
rect -298 778 -245 779
tri -245 778 -244 779 nw
rect -605 771 -546 778
tri -605 766 -600 771 ne
rect -600 766 -546 771
tri -546 766 -534 778 sw
tri -499 766 -487 778 ne
rect -487 766 -259 778
tri -757 764 -755 766 sw
tri -600 764 -598 766 ne
rect -598 764 -534 766
tri -534 764 -532 766 sw
tri -487 764 -485 766 ne
rect -485 764 -259 766
tri -259 764 -245 778 nw
rect -757 730 -755 764
tri -755 730 -721 764 sw
tri -598 762 -596 764 ne
rect -596 762 -532 764
tri -532 762 -530 764 sw
tri -485 762 -483 764 ne
rect -483 762 -291 764
tri -596 730 -564 762 ne
rect -564 732 -530 762
tri -530 732 -500 762 sw
tri -483 732 -453 762 ne
rect -453 732 -291 762
tri -291 732 -259 764 nw
rect -564 730 -500 732
tri -500 730 -498 732 sw
rect -757 722 -721 730
rect -809 718 -721 722
tri -721 718 -709 730 sw
tri -564 718 -552 730 ne
rect -552 728 -498 730
tri -498 728 -496 730 sw
rect -552 718 -496 728
tri -496 718 -486 728 sw
tri -141 718 -131 728 se
rect -131 718 -85 991
tri 7315 970 7336 991 ne
rect 7336 970 7827 991
tri 7827 970 7879 1022 nw
tri 8592 1009 8605 1022 se
rect 8605 1009 8646 1022
tri 8646 1009 8686 1049 nw
tri 8795 1009 8801 1015 se
rect 8801 1009 9720 1015
rect 8035 957 8041 1009
rect 8093 957 8105 1009
rect 8157 970 8607 1009
tri 8607 970 8646 1009 nw
tri 8756 970 8795 1009 se
rect 8795 970 9720 1009
rect 8157 957 8594 970
tri 8594 957 8607 970 nw
tri 8743 957 8756 970 se
rect 8756 969 9720 970
rect 8756 957 8801 969
tri 8735 949 8743 957 se
rect 8743 949 8801 957
tri 8801 949 8821 969 nw
tri 8714 928 8735 949 se
rect 8735 928 8775 949
rect 8628 876 8634 928
rect 8686 876 8698 928
rect 8750 923 8775 928
tri 8775 923 8801 949 nw
rect 8750 876 8756 923
tri 8756 904 8775 923 nw
rect -809 710 -592 718
rect -1224 646 -1222 667
tri -1222 646 -1201 667 sw
rect -757 696 -592 710
tri -592 696 -570 718 sw
tri -552 696 -530 718 ne
rect -530 696 -486 718
tri -486 696 -464 718 sw
tri -163 696 -141 718 se
rect -141 708 -85 718
rect -141 696 -97 708
tri -97 696 -85 708 nw
rect 0 842 11256 848
rect 0 790 7975 842
rect 8027 790 8079 842
rect 8131 836 11256 842
rect 8131 802 8692 836
rect 8726 802 9188 836
rect 9222 802 11256 836
rect 8131 790 11256 802
rect 0 773 11256 790
rect 0 721 7975 773
rect 8027 721 8079 773
rect 8131 764 11256 773
rect 8131 730 8692 764
rect 8726 730 9188 764
rect 9222 730 11256 764
rect 8131 721 11256 730
rect 0 704 11256 721
rect -757 688 -570 696
tri -570 688 -562 696 sw
tri -530 688 -522 696 ne
rect -522 688 -143 696
rect -757 672 -562 688
tri -562 672 -546 688 sw
tri -522 672 -506 688 ne
rect -506 672 -143 688
rect -757 667 -742 672
tri -742 667 -737 672 nw
tri -612 667 -607 672 ne
rect -607 667 -546 672
tri -546 667 -541 672 sw
tri -506 667 -501 672 ne
rect -501 667 -143 672
rect -809 652 -757 658
tri -757 652 -742 667 nw
tri -607 652 -592 667 ne
rect -592 662 -541 667
tri -541 662 -536 667 sw
tri -501 662 -496 667 ne
rect -496 662 -143 667
rect -592 652 -536 662
tri -536 652 -526 662 sw
tri -496 652 -486 662 ne
rect -486 652 -143 662
tri -592 646 -586 652 ne
rect -586 650 -526 652
tri -526 650 -524 652 sw
tri -486 650 -484 652 ne
rect -484 650 -143 652
tri -143 650 -97 696 nw
rect 0 652 7975 704
rect 8027 652 8079 704
rect 8131 652 11256 704
rect -586 646 -524 650
tri -524 646 -520 650 sw
rect 0 646 11256 652
rect -1224 621 -1201 646
tri -1201 621 -1176 646 sw
tri -586 622 -562 646 ne
rect -562 622 -520 646
tri -520 622 -496 646 sw
tri -562 621 -561 622 ne
rect -561 621 -123 622
tri -1224 616 -1219 621 ne
rect -1219 616 -609 621
tri -609 616 -604 621 sw
tri -561 616 -556 621 ne
rect -556 616 -123 621
rect -1359 593 -1302 599
rect -1411 587 -1302 593
tri -1219 592 -1195 616 ne
rect -1195 592 -604 616
tri -604 592 -580 616 sw
tri -556 592 -532 616 ne
rect -532 592 -241 616
tri -1195 587 -1190 592 ne
rect -1190 587 -580 592
tri -623 582 -618 587 ne
rect -618 582 -580 587
tri -580 582 -570 592 sw
tri -532 582 -522 592 ne
rect -522 582 -241 592
rect -207 582 -169 616
rect -135 582 -123 616
rect 9686 612 9849 618
tri -618 578 -614 582 ne
rect -614 578 -570 582
tri -570 578 -566 582 sw
tri -522 578 -518 582 ne
rect -518 578 -123 582
tri 5002 578 5011 587 se
rect 5011 578 5805 587
tri -614 551 -587 578 ne
rect -587 576 -566 578
tri -566 576 -564 578 sw
tri -518 576 -516 578 ne
rect -516 576 -123 578
tri 5000 576 5002 578 se
rect 5002 576 5805 578
rect -587 562 -564 576
tri -564 562 -550 576 sw
tri 4986 562 5000 576 se
rect 5000 562 5805 576
rect -587 551 -550 562
tri -550 551 -539 562 sw
tri 1906 551 1917 562 se
rect 1917 551 1923 562
rect -1593 545 -796 551
rect -1541 537 -1493 545
rect -1441 539 -796 545
tri -587 544 -580 551 ne
rect -580 544 -539 551
tri -539 544 -532 551 sw
tri 1899 544 1906 551 se
rect 1906 544 1923 551
rect -1541 503 -1514 537
rect -1441 505 -1262 539
rect -1228 505 -1138 539
rect -1104 505 -796 539
tri -580 528 -564 544 ne
rect -564 528 1035 544
tri 1035 528 1051 544 sw
tri 1281 528 1297 544 se
rect 1297 528 1923 544
tri -564 510 -546 528 ne
rect -546 510 1923 528
rect 1975 510 1987 562
rect 2039 510 2045 562
tri 4968 544 4986 562 se
rect 4986 544 5805 562
rect -1541 493 -1493 503
rect -1441 493 -796 505
tri 1021 494 1037 510 ne
rect 1037 494 1290 510
tri 1290 494 1306 510 nw
rect -1593 468 -796 493
rect 2878 492 2884 544
rect 2936 492 2948 544
rect 3000 535 5805 544
rect 5857 535 5869 587
rect 5921 535 5927 587
rect 9686 578 9731 612
rect 9765 578 9803 612
rect 9837 578 9849 612
rect 9686 572 9849 578
rect 3000 510 5008 535
tri 5008 510 5033 535 nw
rect 3000 492 3006 510
tri 3006 492 3024 510 nw
rect -1541 459 -1493 468
rect -1441 467 -796 468
rect -1541 425 -1514 459
rect -1441 433 -1262 467
rect -1228 433 -1138 467
rect -1104 433 -796 467
rect -1541 416 -1493 425
rect -1441 416 -796 433
rect -1593 391 -796 416
rect 8172 406 8178 458
rect 8230 406 8242 458
rect 8294 406 8300 458
rect -1541 381 -1493 391
rect -1541 347 -1514 381
rect -1541 339 -1493 347
rect -1441 339 -796 391
rect -1593 336 -796 339
rect -1593 314 -1441 336
rect -1541 304 -1493 314
rect -1541 270 -1514 304
rect -1541 262 -1493 270
rect -1593 237 -1441 262
rect -1541 227 -1493 237
rect -1541 193 -1514 227
rect -1541 185 -1493 193
rect -1593 179 -1441 185
rect -1135 143 -1083 149
rect -1321 90 -1275 102
rect -1321 56 -1315 90
rect -1281 56 -1275 90
rect -1321 18 -1275 56
tri -1083 120 -1067 136 sw
rect 0 120 8127 322
rect 8193 247 8199 299
rect 8251 247 8266 299
rect 8318 247 8332 299
rect 8384 247 8390 299
rect 8193 201 8390 247
rect 8193 149 8199 201
rect 8251 149 8266 201
rect 8318 149 8332 201
rect 8384 149 8390 201
rect -1083 101 -1067 120
tri -1067 101 -1048 120 sw
rect -1083 95 -856 101
rect -1083 91 -974 95
rect -1135 79 -974 91
rect -1083 61 -974 79
rect -940 61 -902 95
rect -868 61 -856 95
rect -1083 55 -856 61
rect 6213 86 6262 92
rect 6314 86 6326 92
rect -1083 52 -1052 55
tri -1052 52 -1049 55 nw
rect 6213 52 6225 86
rect 6259 52 6262 86
rect -1083 40 -1064 52
tri -1064 40 -1052 52 nw
rect 6213 40 6262 52
rect 6314 40 6326 52
rect 6378 40 6384 92
rect 6861 40 7889 92
rect -1135 21 -1083 27
tri -1083 21 -1064 40 nw
rect -1321 -16 -1315 18
rect -1281 -16 -1275 18
rect -1321 -95 -1275 -16
rect -1131 -24 -999 -18
rect -1131 -30 -1051 -24
rect -1131 -64 -1125 -30
rect -1091 -64 -1051 -30
tri -1275 -95 -1255 -75 sw
rect -1131 -76 -1051 -64
rect -1131 -90 -999 -76
tri -1321 -102 -1314 -95 ne
rect -1314 -102 -1255 -95
tri -1255 -102 -1248 -95 sw
rect -1131 -102 -1051 -90
tri -1314 -136 -1280 -102 ne
rect -1280 -136 -1248 -102
tri -1248 -136 -1214 -102 sw
rect -1131 -136 -1125 -102
rect -1091 -136 -1051 -102
tri -1280 -161 -1255 -136 ne
rect -1255 -157 -1214 -136
tri -1214 -157 -1193 -136 sw
rect -1131 -142 -1051 -136
rect -1131 -148 -999 -142
rect -1255 -161 -1193 -157
tri -1193 -161 -1189 -157 sw
tri -1255 -177 -1239 -161 ne
rect -1239 -177 -1189 -161
tri -1189 -177 -1173 -161 sw
tri -1239 -183 -1233 -177 ne
rect -1233 -183 -998 -177
rect -1411 -189 -1359 -183
tri -1233 -202 -1214 -183 ne
rect -1214 -202 -1116 -183
tri -1359 -217 -1344 -202 sw
tri -1214 -217 -1199 -202 ne
rect -1199 -217 -1116 -202
rect -1082 -217 -1044 -183
rect -1010 -217 -998 -183
rect -1359 -233 -1344 -217
tri -1344 -233 -1328 -217 sw
tri -1199 -223 -1193 -217 ne
rect -1193 -223 -998 -217
rect -1359 -241 -1328 -233
rect -1411 -253 -1328 -241
tri -1328 -253 -1308 -233 sw
tri -751 -253 -731 -233 se
rect -731 -253 2680 -233
rect -1359 -285 2680 -253
rect 2732 -285 2744 -233
rect 2796 -285 2802 -233
rect -1359 -305 -729 -285
tri -729 -305 -709 -285 nw
rect -1411 -311 -1354 -305
tri -1354 -311 -1348 -305 nw
tri -1300 -341 -1294 -335 se
rect -1294 -341 -1230 -335
rect -1424 -347 -1230 -341
rect -1424 -381 -1412 -347
rect -1378 -381 -1340 -347
rect -1306 -381 -1230 -347
rect -1424 -387 -1230 -381
rect -1178 -387 -1166 -335
rect -1114 -387 -1108 -335
rect -1135 -579 -933 -539
rect -1360 -604 -877 -598
rect -1360 -638 -1348 -604
rect -1314 -638 -1263 -604
rect -1229 -638 -1178 -604
rect -1144 -638 -1093 -604
rect -1059 -638 -1008 -604
rect -974 -638 -923 -604
rect -889 -638 -877 -604
rect -1360 -644 -877 -638
<< rmetal1 >>
rect 9575 2771 9627 2772
rect 9575 2770 9576 2771
rect 9626 2770 9627 2771
rect 9575 2733 9576 2734
rect 9626 2733 9627 2734
rect 9575 2732 9627 2733
rect 9426 1830 9428 1831
rect 9464 1830 9466 1831
rect 9426 1780 9427 1830
rect 9465 1780 9466 1830
rect 9426 1779 9428 1780
rect 9464 1779 9466 1780
rect 9829 1753 9881 1754
rect 9829 1752 9830 1753
rect 9880 1752 9881 1753
rect 9829 1715 9830 1716
rect 9880 1715 9881 1716
rect 9829 1714 9881 1715
rect 9363 1674 9365 1675
rect 9401 1674 9403 1675
rect 9363 1624 9364 1674
rect 9402 1624 9403 1674
rect 9363 1623 9365 1624
rect 9401 1623 9403 1624
rect 9429 1597 9481 1598
rect 9429 1596 9430 1597
rect 9480 1596 9481 1597
rect 9429 1559 9430 1560
rect 9480 1559 9481 1560
rect 9429 1558 9481 1559
rect 9561 1532 9563 1533
rect 9561 1482 9562 1532
rect 9561 1481 9563 1482
rect 9599 1532 9601 1533
rect 9600 1482 9601 1532
rect 9599 1481 9601 1482
<< via1 >>
rect 8864 3565 8916 3617
rect 8928 3565 8980 3617
rect 4530 3375 4582 3427
rect 4594 3375 4646 3427
rect 8726 3362 8778 3414
rect 8790 3362 8842 3414
rect 9548 3362 9600 3414
rect 9612 3362 9664 3414
rect 9587 3196 9639 3248
rect 9651 3196 9703 3248
rect 3556 3137 3608 3189
rect 3620 3137 3672 3189
rect 4530 3137 4582 3189
rect 4594 3137 4646 3189
rect 8726 3103 8778 3155
rect 8790 3103 8842 3155
rect 11287 3112 11339 3164
rect 6635 3027 6687 3079
rect 6699 3027 6751 3079
rect 11287 3048 11339 3100
rect 9759 2637 9811 2689
rect 9823 2637 9875 2689
rect 9520 2177 9572 2229
rect 9584 2177 9636 2229
rect -945 2035 -893 2087
rect -945 1971 -893 2023
rect -1413 1886 -1361 1892
rect -1413 1852 -1401 1886
rect -1401 1852 -1367 1886
rect -1367 1852 -1361 1886
rect -1413 1840 -1361 1852
rect -1413 1814 -1361 1826
rect -1413 1780 -1401 1814
rect -1401 1780 -1367 1814
rect -1367 1780 -1361 1814
rect -1413 1774 -1361 1780
rect -1135 1835 -1083 1887
rect 5805 2095 5857 2147
rect 5869 2095 5921 2147
rect 7950 2097 8002 2149
rect 8014 2097 8066 2149
rect 9618 2097 9670 2149
rect 9682 2097 9734 2149
rect 9934 2098 9986 2150
rect 9998 2098 10050 2150
rect 10904 2087 10956 2139
rect 8495 2017 8547 2069
rect 8559 2017 8611 2069
rect 10904 2023 10956 2075
rect -141 1928 -89 1980
rect -141 1864 -89 1916
rect -1135 1771 -1083 1823
rect 11492 1855 11544 1907
rect 1947 1672 1999 1724
rect 2011 1672 2063 1724
rect 6711 1656 6763 1708
rect 6775 1656 6827 1708
rect 7497 1678 7549 1730
rect 7875 1704 7927 1756
rect 7939 1704 7991 1756
rect 9514 1779 9566 1831
rect 9578 1779 9630 1831
rect 9759 1779 9811 1831
rect 9823 1779 9875 1831
rect 11492 1791 11544 1843
rect 7497 1614 7549 1666
rect 8634 1623 8686 1675
rect 8698 1623 8750 1675
rect 3556 1531 3608 1583
rect 3620 1531 3672 1583
rect 6810 1471 6862 1523
rect 1172 1403 1224 1455
rect 1236 1403 1288 1455
rect 6037 1401 6089 1453
rect 6101 1401 6153 1453
rect 6810 1407 6862 1459
rect 7283 1401 7335 1453
rect 7347 1401 7399 1453
rect 8726 1401 8778 1453
rect 8790 1401 8842 1453
rect 9040 1441 9092 1453
rect 9040 1407 9049 1441
rect 9049 1407 9083 1441
rect 9083 1407 9092 1441
rect 9040 1401 9092 1407
rect 9104 1441 9156 1453
rect 9104 1407 9121 1441
rect 9121 1407 9155 1441
rect 9155 1407 9156 1441
rect 9104 1401 9156 1407
rect 1172 1089 1224 1141
rect 1236 1089 1288 1141
rect 6037 1089 6089 1141
rect 6101 1089 6153 1141
rect 6262 1073 6314 1125
rect 6326 1073 6378 1125
rect 8942 1119 8994 1171
rect 11287 1138 11339 1190
rect 8942 1055 8994 1107
rect 9677 1064 9729 1116
rect 9741 1064 9793 1116
rect 11287 1074 11339 1126
rect -827 1012 -775 1018
rect -1413 921 -1361 973
rect -1413 857 -1361 909
rect -827 978 -819 1012
rect -819 978 -785 1012
rect -785 978 -775 1012
rect -827 966 -775 978
rect -827 940 -775 952
rect -827 906 -819 940
rect -819 906 -785 940
rect -785 906 -775 940
rect -827 900 -775 906
rect -1411 659 -1359 711
rect -1411 593 -1359 645
rect -1051 785 -999 795
rect -1051 751 -1049 785
rect -1049 751 -1015 785
rect -1015 751 -999 785
rect -1051 743 -999 751
rect -1051 713 -999 731
rect -1051 679 -1049 713
rect -1049 679 -1015 713
rect -1015 679 -999 713
rect -809 722 -757 774
rect 8041 957 8093 1009
rect 8105 957 8157 1009
rect 8634 876 8686 928
rect 8698 876 8750 928
rect -809 658 -757 710
rect 7975 790 8027 842
rect 8079 790 8131 842
rect 7975 721 8027 773
rect 8079 721 8131 773
rect 7975 652 8027 704
rect 8079 652 8131 704
rect -1593 537 -1541 545
rect -1493 537 -1441 545
rect -1593 503 -1586 537
rect -1586 503 -1552 537
rect -1552 503 -1541 537
rect -1493 503 -1480 537
rect -1480 503 -1441 537
rect 1923 510 1975 562
rect 1987 510 2039 562
rect -1593 493 -1541 503
rect -1493 493 -1441 503
rect 2884 492 2936 544
rect 2948 492 3000 544
rect 5805 535 5857 587
rect 5869 535 5921 587
rect -1593 459 -1541 468
rect -1493 459 -1441 468
rect -1593 425 -1586 459
rect -1586 425 -1552 459
rect -1552 425 -1541 459
rect -1493 425 -1480 459
rect -1480 425 -1441 459
rect -1593 416 -1541 425
rect -1493 416 -1441 425
rect 8178 406 8230 458
rect 8242 406 8294 458
rect -1593 381 -1541 391
rect -1493 381 -1441 391
rect -1593 347 -1586 381
rect -1586 347 -1552 381
rect -1552 347 -1541 381
rect -1493 347 -1480 381
rect -1480 347 -1441 381
rect -1593 339 -1541 347
rect -1493 339 -1441 347
rect -1593 304 -1541 314
rect -1493 304 -1441 314
rect -1593 270 -1586 304
rect -1586 270 -1552 304
rect -1552 270 -1541 304
rect -1493 270 -1480 304
rect -1480 270 -1441 304
rect -1593 262 -1541 270
rect -1493 262 -1441 270
rect -1593 227 -1541 237
rect -1493 227 -1441 237
rect -1593 193 -1586 227
rect -1586 193 -1552 227
rect -1552 193 -1541 227
rect -1493 193 -1480 227
rect -1480 193 -1441 227
rect -1593 185 -1541 193
rect -1493 185 -1441 193
rect -1135 91 -1083 143
rect 8199 247 8251 299
rect 8266 247 8318 299
rect 8332 247 8384 299
rect 8199 149 8251 201
rect 8266 149 8318 201
rect 8332 149 8384 201
rect -1135 27 -1083 79
rect 6262 86 6314 92
rect 6326 86 6378 92
rect 6262 52 6297 86
rect 6297 52 6314 86
rect 6326 52 6331 86
rect 6331 52 6378 86
rect 6262 40 6314 52
rect 6326 40 6378 52
rect -1051 -76 -999 -24
rect -1051 -142 -999 -90
rect -1411 -241 -1359 -189
rect -1411 -305 -1359 -253
rect 2680 -285 2732 -233
rect 2744 -285 2796 -233
rect -1230 -387 -1178 -335
rect -1166 -387 -1114 -335
<< metal2 >>
rect 8858 3565 8864 3617
rect 8916 3565 8928 3617
rect 8980 3565 8986 3617
tri 8858 3534 8889 3565 ne
rect 8889 3534 8930 3565
tri 8930 3534 8961 3565 nw
tri 9381 3534 9401 3554 se
rect 9401 3534 9754 3554
tri 9754 3534 9774 3554 sw
rect 4524 3375 4530 3427
rect 4582 3375 4594 3427
rect 4646 3375 4652 3427
tri 4524 3362 4537 3375 ne
rect 4537 3362 4639 3375
tri 4639 3362 4652 3375 nw
rect 8720 3362 8726 3414
rect 8778 3362 8790 3414
rect 8842 3362 8848 3414
tri 4537 3350 4549 3362 ne
rect 4549 3350 4627 3362
tri 4627 3350 4639 3362 nw
tri 8720 3350 8732 3362 ne
rect 8732 3350 8848 3362
tri 4549 3328 4571 3350 ne
tri 4566 3231 4571 3236 se
rect 4571 3231 4627 3350
tri 8732 3286 8796 3350 ne
tri 4549 3214 4566 3231 se
rect 4566 3214 4627 3231
tri 8779 3214 8796 3231 se
rect 8796 3214 8848 3350
tri 4531 3196 4549 3214 se
rect 4549 3196 4627 3214
tri 4627 3196 4645 3214 sw
tri 8761 3196 8779 3214 se
rect 8779 3196 8848 3214
tri 4524 3189 4531 3196 se
rect 4531 3189 4645 3196
tri 4645 3189 4652 3196 sw
rect 3550 3137 3556 3189
rect 3608 3137 3620 3189
rect 3672 3137 3678 3189
rect 4524 3137 4530 3189
rect 4582 3137 4594 3189
rect 4646 3137 4652 3189
tri 8729 3164 8761 3196 se
rect 8761 3164 8848 3196
tri 8720 3155 8729 3164 se
rect 8729 3155 8848 3164
tri 3550 3105 3582 3137 ne
rect 3582 3105 3646 3137
tri 3646 3105 3678 3137 nw
tri 3582 3103 3584 3105 ne
rect 3584 3103 3646 3105
tri 3584 3100 3587 3103 ne
rect 3587 3100 3646 3103
rect 8720 3103 8726 3155
rect 8778 3103 8790 3155
rect 8842 3103 8848 3155
tri 8720 3100 8723 3103 ne
rect 8723 3100 8848 3103
tri 3587 3089 3598 3100 ne
tri -1593 2447 -1511 2529 se
rect -1593 2343 -1511 2447
rect -1593 545 -1441 2343
tri -1441 2279 -1377 2343 nw
rect -945 2087 -893 2093
rect -945 2023 -893 2035
rect -1413 1892 -1361 1898
rect -1413 1826 -1361 1840
rect -1413 973 -1361 1774
rect -1413 909 -1361 921
rect -1413 851 -1361 857
rect -1135 1887 -1083 1893
rect -1135 1823 -1083 1835
rect -1541 493 -1493 545
rect -1593 468 -1441 493
rect -1541 416 -1493 468
rect -1593 391 -1441 416
rect -1541 339 -1493 391
rect -1593 314 -1441 339
rect -1541 262 -1493 314
rect -1593 237 -1441 262
rect -1541 185 -1493 237
rect -1593 179 -1441 185
rect -1411 711 -1359 717
rect -1411 645 -1359 659
rect -1411 -189 -1359 593
rect -1135 143 -1083 1771
rect -945 1294 -893 1971
rect -141 1980 -89 1986
rect -141 1916 -89 1928
rect -141 1809 -89 1864
tri -89 1809 -67 1831 sw
tri -141 1779 -111 1809 ne
rect -111 1779 -67 1809
tri -67 1779 -37 1809 sw
tri -111 1756 -88 1779 ne
rect -88 1756 -37 1779
tri -37 1756 -14 1779 sw
tri -88 1735 -67 1756 ne
rect -67 1746 -14 1756
tri -14 1746 -4 1756 sw
rect -67 1735 -4 1746
tri -67 1730 -62 1735 ne
rect -62 1730 -4 1735
tri -62 1724 -56 1730 ne
rect -56 1660 -4 1730
rect 1941 1672 1947 1724
rect 1999 1672 2011 1724
rect 2063 1672 2069 1724
tri 1941 1660 1953 1672 ne
rect 1953 1660 2046 1672
tri 1953 1656 1957 1660 ne
rect 1957 1656 2046 1660
tri 2046 1656 2062 1672 nw
tri 1957 1643 1970 1656 ne
rect 1166 1403 1172 1455
rect 1224 1403 1236 1455
rect 1288 1403 1294 1455
tri -945 1272 -923 1294 ne
rect -923 1272 -893 1294
tri -893 1272 -849 1316 sw
tri -923 1242 -893 1272 ne
rect -893 1242 -849 1272
tri -893 1198 -849 1242 ne
tri -849 1214 -791 1272 sw
rect -849 1198 -791 1214
tri -791 1198 -775 1214 sw
tri -849 1190 -841 1198 ne
rect -841 1190 -775 1198
tri -841 1176 -827 1190 ne
rect -827 1018 -775 1190
rect 1166 1141 1294 1403
rect 1166 1089 1172 1141
rect 1224 1089 1236 1141
rect 1288 1089 1294 1141
rect -827 952 -775 966
rect -827 894 -775 900
rect -1135 79 -1083 91
rect -1135 21 -1083 27
rect -1051 795 -999 801
rect -1051 731 -999 743
rect -1051 -24 -999 679
rect -812 774 -756 780
rect -812 771 -809 774
rect -757 771 -756 774
rect -812 710 -756 715
rect -812 691 -809 710
rect -757 691 -756 710
rect -812 626 -756 635
tri 1942 587 1970 615 se
rect 1970 587 2033 1656
tri 2033 1643 2046 1656 nw
tri 3582 1615 3598 1631 se
rect 3598 1615 3646 3100
tri 8723 3079 8744 3100 ne
rect 8744 3079 8848 3100
rect 6629 3027 6635 3079
rect 6687 3027 6699 3079
rect 6751 3027 6757 3079
tri 8744 3048 8775 3079 ne
rect 8775 3048 8848 3079
tri 8775 3027 8796 3048 ne
tri 6680 3002 6705 3027 ne
rect 5799 2095 5805 2147
rect 5857 2095 5869 2147
rect 5921 2095 5927 2147
tri 5799 2087 5807 2095 ne
rect 5807 2087 5919 2095
tri 5919 2087 5927 2095 nw
tri 5807 2075 5819 2087 ne
rect 5819 2075 5907 2087
tri 5907 2075 5919 2087 nw
tri 5819 2069 5825 2075 ne
rect 5825 2069 5901 2075
tri 5901 2069 5907 2075 nw
tri 5825 2062 5832 2069 ne
rect 5832 2062 5894 2069
tri 5894 2062 5901 2069 nw
tri 5832 2053 5841 2062 ne
tri 3581 1614 3582 1615 se
rect 3582 1614 3646 1615
tri 3646 1614 3647 1615 sw
tri 3550 1583 3581 1614 se
rect 3581 1583 3647 1614
tri 3647 1583 3678 1614 sw
rect 3550 1531 3556 1583
rect 3608 1531 3620 1583
rect 3672 1531 3678 1583
tri 5832 620 5841 629 se
rect 5841 620 5894 2062
rect 6705 1730 6757 3027
rect 7944 2097 7950 2149
rect 8002 2097 8014 2149
rect 8066 2097 8072 2149
rect 7944 2087 8034 2097
tri 8034 2087 8044 2097 nw
rect 7944 2075 8022 2087
tri 8022 2075 8034 2087 nw
rect 7944 2069 8016 2075
tri 8016 2069 8022 2075 nw
tri 7914 1779 7944 1809 se
rect 7944 1779 7991 2069
tri 7991 2044 8016 2069 nw
rect 8489 2017 8495 2069
rect 8547 2017 8559 2069
rect 8611 2017 8617 2069
rect 8489 1954 8617 2017
rect 8489 1920 8583 1954
tri 8583 1920 8617 1954 nw
tri 8476 1907 8489 1920 se
rect 8489 1907 8570 1920
tri 8570 1907 8583 1920 nw
tri 8424 1855 8476 1907 se
rect 8476 1855 8518 1907
tri 8518 1855 8570 1907 nw
tri 8412 1843 8424 1855 se
rect 8424 1843 8506 1855
tri 8506 1843 8518 1855 nw
tri 8400 1831 8412 1843 se
rect 8412 1831 8494 1843
tri 8494 1831 8506 1843 nw
tri 8395 1826 8400 1831 se
rect 8400 1826 8489 1831
tri 8489 1826 8494 1831 nw
tri 8348 1779 8395 1826 se
rect 8395 1779 8442 1826
tri 8442 1779 8489 1826 nw
tri 7891 1756 7914 1779 se
rect 7914 1756 7991 1779
tri 8331 1762 8348 1779 se
rect 8348 1762 8395 1779
tri 7991 1756 7997 1762 sw
tri 6757 1730 6760 1733 sw
rect 7497 1730 7549 1736
rect 6705 1708 6760 1730
tri 6760 1708 6782 1730 sw
rect 6705 1656 6711 1708
rect 6763 1656 6775 1708
rect 6827 1656 6833 1708
rect 7869 1704 7875 1756
rect 7927 1704 7939 1756
rect 7991 1704 7997 1756
tri 8302 1733 8331 1762 se
rect 8331 1733 8395 1762
tri 8301 1732 8302 1733 se
rect 8302 1732 8395 1733
tri 8395 1732 8442 1779 nw
tri 8277 1708 8301 1732 se
rect 8301 1708 8338 1732
tri 8273 1704 8277 1708 se
rect 8277 1704 8338 1708
rect 7497 1666 7549 1678
tri 8244 1675 8273 1704 se
rect 8273 1675 8338 1704
tri 8338 1675 8395 1732 nw
tri 7496 1608 7497 1609 se
rect 7497 1608 7549 1614
tri 7475 1587 7496 1608 se
rect 7496 1587 7549 1608
tri 7437 1549 7475 1587 se
rect 7475 1549 7511 1587
tri 7511 1549 7549 1587 nw
tri 8233 1664 8244 1675 se
rect 8244 1664 8327 1675
tri 8327 1664 8338 1675 nw
rect 8233 1656 8319 1664
tri 8319 1656 8327 1664 nw
tri 7417 1529 7437 1549 se
rect 7437 1529 7491 1549
tri 7491 1529 7511 1549 nw
rect 6804 1523 6865 1529
rect 6804 1471 6810 1523
rect 6862 1471 6865 1523
tri 7363 1475 7417 1529 se
rect 7417 1475 7437 1529
tri 7437 1475 7491 1529 nw
rect 6804 1459 6865 1471
rect 6031 1401 6037 1453
rect 6089 1401 6101 1453
rect 6153 1401 6159 1453
rect 6031 1141 6159 1401
rect 6804 1407 6810 1459
rect 6862 1407 6865 1459
tri 7341 1453 7363 1475 se
rect 7363 1453 7415 1475
tri 7415 1453 7437 1475 nw
rect 6804 1214 6865 1407
rect 7277 1401 7283 1453
rect 7335 1401 7347 1453
rect 7399 1401 7405 1453
tri 7405 1443 7415 1453 nw
tri 6865 1215 6932 1282 sw
rect 8024 1216 8033 1272
rect 8089 1216 8113 1272
rect 8169 1216 8178 1272
tri 8024 1215 8025 1216 ne
rect 8025 1215 8167 1216
tri 8025 1214 8026 1215 ne
rect 8026 1214 8167 1215
tri 8026 1205 8035 1214 ne
rect 8035 1205 8167 1214
tri 8167 1205 8178 1216 nw
rect 6031 1089 6037 1141
rect 6089 1089 6101 1141
rect 6153 1089 6159 1141
rect 6256 1073 6262 1125
rect 6314 1073 6326 1125
rect 6378 1073 6384 1125
rect 6256 1055 6334 1073
tri 6334 1055 6352 1073 nw
tri 1929 574 1942 587 se
rect 1942 574 2033 587
tri 5799 587 5832 620 se
rect 5832 587 5894 620
tri 5894 587 5927 620 sw
tri 1917 562 1929 574 se
rect 1929 562 2033 574
tri 2033 562 2045 574 sw
rect 1917 510 1923 562
rect 1975 510 1987 562
rect 2039 510 2045 562
rect 2878 492 2884 544
rect 2936 492 2948 544
rect 3000 492 3006 544
rect 5799 535 5805 587
rect 5857 535 5869 587
rect 5921 535 5927 587
tri 2879 458 2913 492 ne
rect 2913 458 2975 492
tri 2975 461 3006 492 nw
tri 2913 449 2922 458 ne
rect -1051 -90 -999 -76
rect -1051 -148 -999 -142
tri 2869 -148 2922 -95 se
rect 2922 -112 2975 458
rect 6256 92 6327 1055
tri 6327 1048 6334 1055 nw
rect 8035 1009 8163 1205
tri 8163 1201 8167 1205 nw
rect 8035 957 8041 1009
rect 8093 957 8105 1009
rect 8157 957 8163 1009
rect 7973 842 8131 848
rect 7973 790 7975 842
rect 8027 790 8079 842
rect 7973 773 8131 790
rect 7973 721 7975 773
rect 8027 721 8079 773
rect 7973 704 8131 721
rect 7973 652 7975 704
rect 8027 652 8079 704
rect 7973 303 8131 652
tri 8208 458 8233 483 se
rect 8233 458 8300 1656
tri 8300 1637 8319 1656 nw
rect 8628 1623 8634 1675
rect 8686 1623 8698 1675
rect 8750 1623 8756 1675
rect 8628 928 8692 1623
tri 8692 1598 8717 1623 nw
tri 8771 1453 8796 1478 se
rect 8796 1453 8848 3048
rect 8720 1401 8726 1453
rect 8778 1401 8790 1453
rect 8842 1401 8848 1453
tri 8875 1379 8889 1393 se
rect 8889 1379 8929 3534
tri 8929 3533 8930 3534 nw
tri 9380 3533 9381 3534 se
rect 9381 3533 9774 3534
tri 9774 3533 9775 3534 sw
tri 9366 3519 9380 3533 se
rect 9380 3519 9775 3533
tri 9775 3519 9789 3533 sw
tri 9346 3499 9366 3519 se
rect 9366 3510 9789 3519
rect 9366 3499 9408 3510
tri 9408 3499 9419 3510 nw
tri 9736 3499 9747 3510 ne
rect 9747 3499 9789 3510
rect 9346 3362 9390 3499
tri 9390 3481 9408 3499 nw
tri 9747 3481 9765 3499 ne
rect 9765 3481 9789 3499
tri 9765 3457 9789 3481 ne
tri 9789 3457 9851 3519 sw
rect 9789 3414 9851 3457
tri 9851 3414 9894 3457 sw
tri 9390 3362 9422 3394 sw
rect 9542 3362 9548 3414
rect 9600 3362 9612 3414
rect 9664 3362 9670 3414
rect 9789 3413 9894 3414
tri 9894 3413 9895 3414 sw
rect 9346 3332 9422 3362
tri 9422 3332 9452 3362 sw
tri 9574 3332 9604 3362 ne
rect 9346 3319 9495 3332
tri 9346 3287 9378 3319 ne
rect 9378 3287 9495 3319
tri 9456 3271 9472 3287 ne
rect 9472 3271 9495 3287
tri 9472 3248 9495 3271 ne
tri 9581 3248 9604 3271 se
rect 9604 3248 9670 3362
tri 9670 3248 9709 3287 sw
rect 9581 3196 9587 3248
rect 9639 3196 9651 3248
rect 9703 3196 9709 3248
rect 11287 3164 11339 3178
rect 11287 3100 11339 3112
tri 9616 2703 9682 2769 se
rect 9682 2717 9755 2769
tri 9682 2703 9696 2717 nw
tri 9602 2689 9616 2703 se
rect 9616 2689 9668 2703
tri 9668 2689 9682 2703 nw
tri 9588 2675 9602 2689 se
rect 9602 2675 9654 2689
tri 9654 2675 9668 2689 nw
tri 9552 2507 9588 2543 se
rect 9588 2507 9634 2675
tri 9634 2655 9654 2675 nw
rect 9753 2637 9759 2689
rect 9811 2637 9823 2689
rect 9875 2637 9881 2689
tri 9804 2612 9829 2637 ne
rect 9468 2451 9477 2507
rect 9533 2451 9557 2507
rect 9613 2451 9634 2507
rect 9514 2177 9520 2229
rect 9572 2177 9584 2229
rect 9636 2177 9642 2229
tri 9514 2169 9522 2177 ne
rect 9522 2023 9574 2177
tri 9574 2151 9600 2177 nw
rect 9612 2097 9618 2149
rect 9670 2097 9682 2149
rect 9734 2097 9740 2149
tri 9642 2087 9652 2097 ne
rect 9652 2087 9740 2097
tri 9652 2075 9664 2087 ne
rect 9664 2075 9740 2087
tri 9664 2068 9671 2075 ne
rect 9671 2067 9740 2075
tri 9574 2023 9580 2029 sw
rect 9522 2007 9580 2023
tri 9522 1967 9562 2007 ne
rect 9562 1967 9580 2007
tri 9580 1967 9636 2023 sw
tri 9562 1955 9574 1967 ne
rect 9574 1955 9636 1967
tri 9574 1945 9584 1955 ne
tri 9583 1855 9584 1856 se
rect 9584 1855 9636 1955
tri 9571 1843 9583 1855 se
rect 9583 1843 9636 1855
tri 9559 1831 9571 1843 se
rect 9571 1831 9636 1843
rect 9508 1779 9514 1831
rect 9566 1779 9578 1831
rect 9630 1779 9636 1831
tri 9029 1420 9034 1425 se
rect 9034 1420 9040 1453
tri 9010 1401 9029 1420 se
rect 9029 1401 9040 1420
rect 9092 1401 9104 1453
rect 9156 1401 9162 1453
tri 8988 1379 9010 1401 se
rect 9010 1379 9062 1401
tri 9062 1379 9084 1401 nw
tri 8831 1335 8875 1379 se
rect 8875 1375 8929 1379
rect 8875 1335 8889 1375
tri 8889 1335 8929 1375 nw
tri 8944 1335 8988 1379 se
rect 8988 1335 9016 1379
tri 8790 1294 8831 1335 se
rect 8831 1294 8848 1335
tri 8848 1294 8889 1335 nw
tri 8942 1333 8944 1335 se
rect 8944 1333 9016 1335
tri 9016 1333 9062 1379 nw
rect 8790 1055 8830 1294
tri 8830 1276 8848 1294 nw
rect 8942 1171 8994 1333
tri 8994 1311 9016 1333 nw
rect 8942 1107 8994 1119
tri 8830 1055 8832 1057 sw
rect 9671 1190 9723 2067
tri 9723 2050 9740 2067 nw
tri 9828 1855 9829 1856 se
rect 9829 1855 9881 2637
tri 9932 2154 10000 2222 se
rect 10000 2154 10052 2724
rect 10453 2184 10501 2236
tri 9928 2150 9932 2154 se
rect 9932 2150 10052 2154
tri 10052 2150 10056 2154 sw
rect 9928 2098 9934 2150
rect 9986 2098 9998 2150
rect 10050 2098 10056 2150
rect 10904 2139 10956 2145
tri 9816 1843 9828 1855 se
rect 9828 1843 9881 1855
rect 10904 2075 10956 2087
rect 10904 1855 10956 2023
tri 10956 1855 10985 1884 sw
tri 10893 1843 10904 1854 se
rect 10904 1843 10985 1855
tri 10985 1843 10997 1855 sw
tri 9804 1831 9816 1843 se
rect 9816 1831 9881 1843
tri 10881 1831 10893 1843 se
rect 10893 1831 10997 1843
tri 10997 1831 11009 1843 sw
rect 9753 1779 9759 1831
rect 9811 1779 9823 1831
rect 9875 1779 9881 1831
rect 9962 1779 10020 1828
tri 9723 1190 9725 1192 sw
rect 11287 1190 11339 3048
rect 11492 1907 11544 1913
rect 11492 1843 11544 1855
rect 11492 1785 11544 1791
rect 9671 1138 9725 1190
tri 9725 1138 9777 1190 sw
rect 9671 1126 9777 1138
tri 9777 1126 9789 1138 sw
rect 11287 1126 11339 1138
rect 9671 1116 9789 1126
tri 9789 1116 9799 1126 sw
rect 9671 1064 9677 1116
rect 9729 1064 9741 1116
rect 9793 1064 9799 1116
rect 11287 1068 11339 1074
rect 8790 1049 8832 1055
tri 8832 1049 8838 1055 sw
rect 8942 1049 8994 1055
rect 8790 1039 8838 1049
tri 8838 1039 8848 1049 sw
tri 8790 981 8848 1039 ne
tri 8848 1023 8864 1039 sw
rect 8848 981 8864 1023
tri 8864 981 8906 1023 sw
tri 8848 965 8864 981 ne
rect 8864 965 8906 981
tri 8906 965 8922 981 sw
rect 8864 953 8922 965
tri 8922 953 8934 965 sw
tri 8692 928 8717 953 sw
rect 8864 932 8934 953
tri 8934 932 8955 953 sw
rect 8628 876 8634 928
rect 8686 876 8698 928
rect 8750 876 8756 928
rect 8172 406 8178 458
rect 8230 406 8242 458
rect 8294 406 8300 458
tri 8131 303 8184 356 sw
rect 7973 299 8392 303
rect 7973 247 8199 299
rect 8251 247 8266 299
rect 8318 247 8332 299
rect 8384 247 8392 299
rect 7973 244 8392 247
tri 7973 201 8016 244 ne
rect 8016 201 8392 244
tri 8016 149 8068 201 ne
rect 8068 149 8199 201
rect 8251 149 8266 201
rect 8318 149 8332 201
rect 8384 149 8392 201
tri 8068 145 8072 149 ne
rect 8072 145 8392 149
tri 6327 92 6352 117 sw
rect 6256 40 6262 92
rect 6314 40 6326 92
rect 6378 40 6384 92
tri 2852 -165 2869 -148 se
rect 2869 -165 2922 -148
tri 2922 -165 2975 -112 nw
tri 2784 -233 2852 -165 se
rect 2852 -233 2854 -165
tri 2854 -233 2922 -165 nw
rect -1411 -253 -1359 -241
rect -1411 -311 -1359 -305
rect -1215 -272 -1159 -263
tri -1236 -335 -1215 -314 se
rect 2674 -285 2680 -233
rect 2732 -285 2744 -233
rect 2796 -285 2802 -233
tri 2802 -285 2854 -233 nw
rect -1215 -335 -1159 -328
tri -1159 -335 -1129 -305 sw
rect -1236 -387 -1230 -335
rect -1178 -352 -1166 -335
rect -1114 -387 -1108 -335
tri -1236 -408 -1215 -387 ne
rect -1215 -417 -1159 -408
tri -1159 -417 -1129 -387 nw
<< via2 >>
rect -812 722 -809 771
rect -809 722 -757 771
rect -757 722 -756 771
rect -812 715 -756 722
rect -812 658 -809 691
rect -809 658 -757 691
rect -757 658 -756 691
rect -812 635 -756 658
rect 8033 1216 8089 1272
rect 8113 1216 8169 1272
rect 9477 2451 9533 2507
rect 9557 2451 9613 2507
rect -1215 -328 -1159 -272
rect -1215 -387 -1178 -352
rect -1178 -387 -1166 -352
rect -1166 -387 -1159 -352
rect -1215 -408 -1159 -387
<< metal3 >>
rect 9472 2507 9618 2512
rect 9472 2506 9477 2507
rect 9533 2506 9557 2507
rect -907 2442 -901 2506
rect -837 2442 -821 2506
rect -757 2442 -751 2506
rect 9462 2442 9468 2506
rect 9533 2451 9548 2506
rect 9613 2451 9618 2507
rect 9532 2442 9548 2451
rect 9612 2442 9618 2451
tri -907 2352 -817 2442 ne
rect -1258 1211 -1252 1275
rect -1188 1211 -1172 1275
rect -1108 1211 -1102 1275
tri -1258 1173 -1220 1211 ne
rect -1220 1173 -1140 1211
tri -1140 1173 -1102 1211 nw
rect -1220 -272 -1154 1173
tri -1154 1159 -1140 1173 nw
rect -817 771 -751 2442
rect 8012 1275 8174 1277
rect 8012 1211 8023 1275
rect 8087 1272 8103 1275
rect 8167 1272 8174 1275
rect 8089 1216 8103 1272
rect 8169 1216 8174 1272
rect 8087 1211 8103 1216
rect 8167 1211 8174 1216
rect -817 715 -812 771
rect -756 715 -751 771
rect -817 691 -751 715
rect -817 635 -812 691
rect -756 635 -751 691
rect -817 630 -751 635
rect -1220 -328 -1215 -272
rect -1159 -328 -1154 -272
rect -1220 -352 -1154 -328
rect -1220 -408 -1215 -352
rect -1159 -408 -1154 -352
rect -1220 -413 -1154 -408
<< via3 >>
rect -901 2442 -837 2506
rect -821 2442 -757 2506
rect 9468 2451 9477 2506
rect 9477 2451 9532 2506
rect 9548 2451 9557 2506
rect 9557 2451 9612 2506
rect 9468 2442 9532 2451
rect 9548 2442 9612 2451
rect -1252 1211 -1188 1275
rect -1172 1211 -1108 1275
rect 8023 1272 8087 1275
rect 8103 1272 8167 1275
rect 8023 1216 8033 1272
rect 8033 1216 8087 1272
rect 8103 1216 8113 1272
rect 8113 1216 8167 1272
rect 8023 1211 8087 1216
rect 8103 1211 8167 1216
<< metal4 >>
rect -902 2506 9613 2507
rect -902 2442 -901 2506
rect -837 2442 -821 2506
rect -757 2442 9468 2506
rect 9532 2442 9548 2506
rect 9612 2442 9613 2506
rect -902 2441 9613 2442
rect -1305 1275 8168 1276
rect -1305 1211 -1252 1275
rect -1188 1211 -1172 1275
rect -1108 1211 8023 1275
rect 8087 1211 8103 1275
rect 8167 1211 8168 1275
rect -1305 1210 8168 1211
use sky130_fd_io__com_pdpredrvr_pbiasv2  sky130_fd_io__com_pdpredrvr_pbiasv2_0
timestamp 1663361622
transform -1 0 20068 0 1 -2980
box 11364 2930 20068 5671
use sky130_fd_io__gpiov2_octl_mux  sky130_fd_io__gpiov2_octl_mux_0
timestamp 1663361622
transform 1 0 -1627 0 -1 3513
box 1191 1040 1945 3147
use sky130_fd_io__gpiov2_pdpredrvr_strong_nr2  sky130_fd_io__gpiov2_pdpredrvr_strong_nr2_0
timestamp 1663361622
transform 1 0 3465 0 -1 -331
box 4658 -2162 7919 -248
use sky130_fd_io__gpiov2_pdpredrvr_strong_nr3  sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0
timestamp 1663361622
transform -1 0 12458 0 1 3202
box 1018 -1305 3472 722
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1663361622
transform -1 0 -1117 0 -1 418
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1663361622
transform -1 0 -1117 0 -1 2582
box -46 24 399 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1663361622
transform 1 0 -1299 0 -1 418
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1663361622
transform 1 0 -1299 0 -1 2582
box -42 24 569 1116
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1663361622
transform 0 1 9429 1 0 1506
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1663361622
transform 0 1 9829 -1 0 1806
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_2
timestamp 1663361622
transform 1 0 9509 0 1 1481
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1663361622
transform -1 0 9455 0 -1 1675
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1663361622
transform 0 -1 9627 1 0 2680
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_2
timestamp 1663361622
transform -1 0 9518 0 1 1779
box 0 0 1 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808139  sky130_fd_pr__model__nfet_highvoltage__example_55959141808139_0
timestamp 1663361622
transform 1 0 8867 0 1 1623
box -15 0 311 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808183  sky130_fd_pr__model__nfet_highvoltage__example_55959141808183_0
timestamp 1663361622
transform 1 0 9247 0 1 1623
box -15 0 121 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808369  sky130_fd_pr__model__nfet_highvoltage__example_55959141808369_0
timestamp 1663361622
transform 1 0 -1093 0 -1 596
box -1 0 121 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808643  sky130_fd_pr__model__nfet_highvoltage__example_55959141808643_0
timestamp 1663361622
transform 1 0 -1373 0 -1 540
box -1 0 101 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_0
timestamp 1663361622
transform 1 0 8867 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_1
timestamp 1663361622
transform -1 0 9163 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808184  sky130_fd_pr__model__pfet_highvoltage__example_55959141808184_0
timestamp 1663361622
transform 1 0 9247 0 -1 1363
box -15 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808371  sky130_fd_pr__model__pfet_highvoltage__example_55959141808371_0
timestamp 1663361622
transform 1 0 -1093 0 -1 994
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808371  sky130_fd_pr__model__pfet_highvoltage__example_55959141808371_1
timestamp 1663361622
transform 1 0 -1093 0 1 1062
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808642  sky130_fd_pr__model__pfet_highvoltage__example_55959141808642_0
timestamp 1663361622
transform 1 0 -1373 0 -1 1394
box -1 0 101 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1663361622
transform 0 -1 -1228 -1 0 539
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1663361622
transform 0 -1 -1104 -1 0 539
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1663361622
transform 0 -1 -1104 1 0 1184
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1663361622
transform 0 -1 9222 -1 0 836
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1663361622
transform 1 0 9049 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1663361622
transform 1 0 8876 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1663361622
transform 0 1 9188 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1663361622
transform 0 1 8808 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1663361622
transform 1 0 8781 0 -1 1209
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1663361622
transform 1 0 6225 0 1 52
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1663361622
transform 1 0 9363 0 -1 1523
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1663361622
transform 0 -1 8726 -1 0 836
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1663361622
transform 1 0 9508 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1663361622
transform -1 0 9881 0 1 2637
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1663361622
transform -1 0 9881 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1663361622
transform -1 0 8848 0 1 1401
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1663361622
transform 1 0 6256 0 1 40
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1663361622
transform 1 0 6256 0 1 1073
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1663361622
transform 1 0 8172 0 1 406
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1663361622
transform 1 0 8628 0 1 876
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1663361622
transform 1 0 8628 0 1 1623
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1663361622
transform 1 0 6629 0 1 3027
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1663361622
transform 1 0 6705 0 1 1656
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1663361622
transform 0 -1 -999 -1 0 762
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1663361622
transform 0 1 8894 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1663361622
transform 0 1 9070 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1663361622
transform 0 1 9247 1 0 1395
box 0 0 1 1
<< labels >>
flabel metal2 s 10453 2184 10501 2236 7 FreeSans 300 180 0 0 PD_H[3]
port 1 nsew
flabel metal2 s 9962 1779 10020 1828 7 FreeSans 300 180 0 0 PD_H[2]
port 2 nsew
flabel metal1 s 11216 2271 11256 2473 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 11216 2797 11256 2999 7 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 7286 3511 7326 3657 7 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 11235 2372 11235 2372 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 11216 646 11256 848 7 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 8087 120 8127 322 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 11216 1243 11256 1373 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 11216 1859 11256 1989 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 6955 40 7000 92 8 FreeSans 300 180 0 0 DRVLO_H_N
port 5 nsew
flabel metal1 s -964 2185 -918 2231 7 FreeSans 300 180 0 0 SLOW_H
port 6 nsew
flabel metal1 s 8796 1407 8848 1453 6 FreeSans 300 180 0 0 PDEN_H_N
port 7 nsew
flabel metal1 s 0 2271 40 2473 3 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 0 1859 40 1989 3 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 272 1243 312 1373 3 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 0 646 40 848 3 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 0 120 40 322 3 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 0 2797 40 2999 3 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 0 3511 40 3657 7 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s -1047 679 -1015 750 3 FreeSans 520 0 0 0 I2C_MODE_H_N
port 8 nsew
flabel metal1 s -1279 336 -960 394 3 FreeSans 520 0 0 0 VGND
port 9 nsew
flabel metal1 s 10929 1788 10977 1820 3 FreeSans 520 0 0 0 PD_H[4]
port 10 nsew
flabel metal1 s -1135 1251 -933 1291 3 FreeSans 300 90 0 0 VCC_IO
port 4 nsew
flabel metal1 s -1135 1574 -933 1614 3 FreeSans 300 90 0 0 VCC_IO
port 4 nsew
flabel metal1 s -1222 2437 -1151 2488 3 FreeSans 520 0 0 0 VGND
port 9 nsew
flabel metal1 s -1135 -579 -933 -539 3 FreeSans 300 90 0 0 VCC_IO
port 4 nsew
flabel comment s 8277 742 8277 742 0 FreeSans 300 0 0 0 VCC_IO
flabel comment s 8253 210 8253 210 0 FreeSans 300 0 0 0 VGND_IO
flabel comment s 7705 3061 7705 3061 0 FreeSans 300 0 0 0 PDEN_H_N
flabel comment s 8813 3706 8813 3706 0 FreeSans 300 90 0 0 PDEN_H_N
flabel comment s 8812 2082 8812 2082 0 FreeSans 300 90 0 0 PDEN_H_N
flabel comment s 8698 1667 8698 1667 0 FreeSans 300 0 0 0 PBIAS
flabel comment s 6897 1611 6897 1611 0 FreeSans 300 0 0 0 EN_FAST_H_N
flabel comment s 9463 1511 9463 1511 0 FreeSans 300 0 0 0 EN_FAST_H_N
flabel comment s 8310 1126 8310 1126 0 FreeSans 300 0 0 0 EN_FAST_H
flabel comment s 6333 1097 6333 1097 0 FreeSans 300 0 0 0 EN_FAST_H
flabel comment s 9956 1467 9956 1467 0 FreeSans 300 0 0 0 PBIAS
flabel comment s 9841 2135 9841 2135 0 FreeSans 300 90 0 0 EN_FAST2_N0
flabel comment s 9565 1662 9565 1662 0 FreeSans 300 0 0 0 EN_FAST_N1
flabel comment s 9600 2130 9600 2130 0 FreeSans 300 90 0 0 EN_FAST2_N1
<< properties >>
string GDS_END 49061400
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 49012710
<< end >>
