magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 5 0 6 4 C0
port 1 nsew
rlabel  s 0 5 5 5 6 C0
port 1 nsew
rlabel  s 0 4 0 5 4 C0
port 1 nsew
rlabel  s 0 4 5 4 6 C0
port 1 nsew
rlabel  s 0 3 0 4 4 C0
port 1 nsew
rlabel  s 0 2 5 3 6 C0
port 1 nsew
rlabel  s 0 2 0 2 4 C0
port 1 nsew
rlabel  s 0 1 5 2 6 C0
port 1 nsew
rlabel  s 0 0 0 1 2 C0
port 1 nsew
rlabel  s 0 0 6 0 8 C0
port 1 nsew
rlabel  s 5 5 6 5 6 C1
port 2 nsew
rlabel  s 5 3 6 4 6 C1
port 2 nsew
rlabel  s 5 2 6 3 6 C1
port 2 nsew
rlabel  s 5 1 6 2 6 C1
port 2 nsew
rlabel  s 1 5 6 6 6 C1
port 2 nsew
rlabel  s 1 4 6 5 6 C1
port 2 nsew
rlabel  s 1 3 6 3 6 C1
port 2 nsew
rlabel  s 1 2 6 2 6 C1
port 2 nsew
rlabel  s 1 1 6 1 6 C1
port 2 nsew
rlabel metal_blue s 3 4 3 4 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 6 6
string LEFview TRUE
<< end >>
