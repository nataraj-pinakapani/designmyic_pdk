magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 5 6 8 6 DRAIN
port 1 nsew
rlabel  s 2 9 5 9 6 GATE
port 2 nsew
rlabel  s 2 3 5 3 6 GATE
port 2 nsew
rlabel  s 0 10 6 13 6 SOURCE
port 3 nsew
rlabel  s 0 0 6 3 6 SOURCE
port 3 nsew
rlabel rotate s 1 9 1 9 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 8 1 8 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 8 1 8 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 7 1 8 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 7 1 7 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 7 1 7 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 6 1 7 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 6 1 6 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 6 1 6 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 5 1 5 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 5 1 5 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 5 1 5 6 SUBSTRATE
port 4 nsew
rlabel rotate s 1 4 1 4 6 SUBSTRATE
port 4 nsew
rlabel  s 1 4 1 9 6 SUBSTRATE
port 4 nsew
rlabel  s 1 4 1 9 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 6 13
string LEFview TRUE
<< end >>
