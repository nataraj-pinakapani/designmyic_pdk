magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1906 203
rect 30 -17 64 21
<< locali >>
rect 17 337 72 493
rect 203 337 239 493
rect 369 337 407 493
rect 537 337 575 493
rect 705 337 743 493
rect 914 337 952 493
rect 1082 337 1120 493
rect 1257 337 1296 420
rect 1409 337 1478 344
rect 17 303 1478 337
rect 17 163 75 303
rect 109 215 351 269
rect 388 215 710 269
rect 763 215 1091 269
rect 1222 215 1465 269
rect 1564 215 1915 268
rect 17 129 337 163
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 106 371 169 527
rect 278 371 335 527
rect 441 371 503 527
rect 609 371 671 527
rect 815 371 880 527
rect 986 371 1044 527
rect 1157 454 1401 493
rect 1157 371 1223 454
rect 1341 412 1401 454
rect 1511 446 1577 527
rect 1611 412 1647 493
rect 1341 378 1647 412
rect 1609 337 1647 378
rect 1682 371 1744 527
rect 1778 337 1816 493
rect 1609 303 1816 337
rect 1853 307 1915 527
rect 371 123 757 165
rect 795 131 1888 181
rect 371 95 405 123
rect 19 57 405 95
rect 439 51 1113 89
rect 1220 17 1286 97
rect 1392 17 1458 97
rect 1565 17 1631 97
rect 1733 17 1799 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 1564 215 1915 268 6 A1
port 1 nsew signal input
rlabel locali s 1222 215 1465 269 6 A2
port 2 nsew signal input
rlabel locali s 763 215 1091 269 6 B1
port 3 nsew signal input
rlabel locali s 388 215 710 269 6 C1
port 4 nsew signal input
rlabel locali s 109 215 351 269 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1906 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 17 129 337 163 6 Y
port 10 nsew signal output
rlabel locali s 17 163 75 303 6 Y
port 10 nsew signal output
rlabel locali s 17 303 1478 337 6 Y
port 10 nsew signal output
rlabel locali s 1409 337 1478 344 6 Y
port 10 nsew signal output
rlabel locali s 1257 337 1296 420 6 Y
port 10 nsew signal output
rlabel locali s 1082 337 1120 493 6 Y
port 10 nsew signal output
rlabel locali s 914 337 952 493 6 Y
port 10 nsew signal output
rlabel locali s 705 337 743 493 6 Y
port 10 nsew signal output
rlabel locali s 537 337 575 493 6 Y
port 10 nsew signal output
rlabel locali s 369 337 407 493 6 Y
port 10 nsew signal output
rlabel locali s 203 337 239 493 6 Y
port 10 nsew signal output
rlabel locali s 17 337 72 493 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1932 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 976088
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 960678
<< end >>
