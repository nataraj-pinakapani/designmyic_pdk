magic
tech minimum
timestamp 1644097873
<< properties >>
string gencell sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1
string parameter m=1
string library sky130
<< end >>
