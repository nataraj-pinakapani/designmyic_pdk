magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< obsli1 >>
rect 126 1732 1598 1798
rect 126 192 192 1732
rect 528 1330 1196 1396
rect 528 594 594 1330
rect 761 759 963 1165
rect 1130 594 1196 1330
rect 528 528 1196 594
rect 1532 192 1598 1732
rect 126 126 1598 192
<< obsm1 >>
rect 130 1736 1594 1794
rect 130 188 188 1736
rect 532 1334 1192 1392
rect 532 590 590 1334
rect 761 789 963 1135
rect 1134 590 1192 1334
rect 532 532 1192 590
rect 1536 188 1594 1736
rect 130 130 1594 188
<< properties >>
string FIXED_BBOX 0 0 1724 1924
string LEFclass BLOCK
string LEFview TRUE
string gencell sky130_fd_pr__rf_npn_05v5_W1p00L2p00
string library sky130
string parameter m=1
string GDS_END 8763626
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 8739358
<< end >>
