magic
tech sky130B
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_0
timestamp 1663361622
transform -1 0 -165 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_1
timestamp 1663361622
transform 1 0 471 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_2
timestamp 1663361622
transform 1 0 1307 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_3
timestamp 1663361622
transform 1 0 2143 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_4
timestamp 1663361622
transform 1 0 2979 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_5
timestamp 1663361622
transform 1 0 3815 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_6
timestamp 1663361622
transform 1 0 4651 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_7
timestamp 1663361622
transform 1 0 5487 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_8
timestamp 1663361622
transform 1 0 6323 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_9
timestamp 1663361622
transform 1 0 7159 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_10
timestamp 1663361622
transform 1 0 7995 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 8150934
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 8140328
<< end >>
