magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 891 203
rect 30 -17 64 21
<< locali >>
rect 283 325 333 425
rect 563 325 613 425
rect 283 289 613 325
rect 40 215 197 257
rect 231 215 385 255
rect 419 181 468 289
rect 511 215 645 255
rect 679 215 833 257
rect 107 145 468 181
rect 107 129 173 145
rect 275 129 341 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 30 325 81 493
rect 115 359 165 527
rect 199 459 417 493
rect 199 325 249 459
rect 30 291 249 325
rect 367 359 417 459
rect 479 459 697 493
rect 479 359 529 459
rect 647 325 697 459
rect 731 359 781 527
rect 815 325 866 493
rect 647 291 866 325
rect 18 95 73 181
rect 502 145 873 181
rect 502 95 536 145
rect 18 61 536 95
rect 571 17 605 111
rect 639 51 705 145
rect 739 17 773 111
rect 807 51 873 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 679 215 833 257 6 A1
port 1 nsew signal input
rlabel locali s 511 215 645 255 6 A2
port 2 nsew signal input
rlabel locali s 40 215 197 257 6 B1
port 3 nsew signal input
rlabel locali s 231 215 385 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 891 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 275 129 341 145 6 Y
port 9 nsew signal output
rlabel locali s 107 129 173 145 6 Y
port 9 nsew signal output
rlabel locali s 107 145 468 181 6 Y
port 9 nsew signal output
rlabel locali s 419 181 468 289 6 Y
port 9 nsew signal output
rlabel locali s 283 289 613 325 6 Y
port 9 nsew signal output
rlabel locali s 563 325 613 425 6 Y
port 9 nsew signal output
rlabel locali s 283 325 333 425 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1388056
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1380180
<< end >>
