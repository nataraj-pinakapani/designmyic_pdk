magic
tech minimum
timestamp 1644097874
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 5 8
string LEFview TRUE
<< end >>
