magic
tech sky130B
timestamp 1663361622
<< metal4 >>
rect -270 7258 6270 7270
rect -270 7140 -258 7258
rect -140 7140 -19 7258
rect 99 7140 141 7258
rect 259 7140 301 7258
rect 419 7140 461 7258
rect 579 7140 621 7258
rect 739 7140 781 7258
rect 899 7140 941 7258
rect 1059 7140 1101 7258
rect 1219 7140 1261 7258
rect 1379 7140 1421 7258
rect 1539 7140 1581 7258
rect 1699 7140 1741 7258
rect 1859 7140 1901 7258
rect 2019 7140 2061 7258
rect 2179 7140 2221 7258
rect 2339 7140 2381 7258
rect 2499 7140 2541 7258
rect 2659 7140 2701 7258
rect 2819 7140 2861 7258
rect 2979 7140 3021 7258
rect 3139 7140 3181 7258
rect 3299 7140 3341 7258
rect 3459 7140 3501 7258
rect 3619 7140 3661 7258
rect 3779 7140 3821 7258
rect 3939 7140 3981 7258
rect 4099 7140 4141 7258
rect 4259 7140 4301 7258
rect 4419 7140 4461 7258
rect 4579 7140 4621 7258
rect 4739 7140 4781 7258
rect 4899 7140 4941 7258
rect 5059 7140 5101 7258
rect 5219 7140 5261 7258
rect 5379 7140 5421 7258
rect 5539 7140 5581 7258
rect 5699 7140 5741 7258
rect 5859 7140 5901 7258
rect 6019 7140 6140 7258
rect 6258 7140 6270 7258
rect -270 7079 6270 7140
rect -270 6961 -258 7079
rect -140 7000 6140 7079
rect -140 6961 0 7000
rect -270 6919 0 6961
rect -270 6801 -258 6919
rect -140 6801 0 6919
rect -270 6759 0 6801
rect -270 6641 -258 6759
rect -140 6641 0 6759
rect -270 6599 0 6641
rect -270 6481 -258 6599
rect -140 6481 0 6599
rect -270 6439 0 6481
rect -270 6321 -258 6439
rect -140 6321 0 6439
rect -270 6279 0 6321
rect -270 6161 -258 6279
rect -140 6161 0 6279
rect -270 6119 0 6161
rect -270 6001 -258 6119
rect -140 6001 0 6119
rect -270 5959 0 6001
rect -270 5841 -258 5959
rect -140 5841 0 5959
rect -270 5799 0 5841
rect -270 5681 -258 5799
rect -140 5681 0 5799
rect -270 5639 0 5681
rect -270 5521 -258 5639
rect -140 5521 0 5639
rect -270 5479 0 5521
rect -270 5361 -258 5479
rect -140 5361 0 5479
rect -270 5319 0 5361
rect -270 5201 -258 5319
rect -140 5201 0 5319
rect -270 5159 0 5201
rect -270 5041 -258 5159
rect -140 5041 0 5159
rect -270 4999 0 5041
rect -270 4881 -258 4999
rect -140 4881 0 4999
rect -270 4839 0 4881
rect -270 4721 -258 4839
rect -140 4721 0 4839
rect -270 4679 0 4721
rect -270 4561 -258 4679
rect -140 4561 0 4679
rect -270 4519 0 4561
rect -270 4401 -258 4519
rect -140 4401 0 4519
rect -270 4359 0 4401
rect -270 4241 -258 4359
rect -140 4241 0 4359
rect -270 4199 0 4241
rect -270 4081 -258 4199
rect -140 4081 0 4199
rect -270 4039 0 4081
rect -270 3921 -258 4039
rect -140 3921 0 4039
rect -270 3879 0 3921
rect -270 3761 -258 3879
rect -140 3761 0 3879
rect -270 3719 0 3761
rect -270 3601 -258 3719
rect -140 3601 0 3719
rect -270 3559 0 3601
rect -270 3441 -258 3559
rect -140 3441 0 3559
rect -270 3399 0 3441
rect -270 3281 -258 3399
rect -140 3281 0 3399
rect -270 3239 0 3281
rect -270 3121 -258 3239
rect -140 3121 0 3239
rect -270 3079 0 3121
rect -270 2961 -258 3079
rect -140 2961 0 3079
rect -270 2919 0 2961
rect -270 2801 -258 2919
rect -140 2801 0 2919
rect -270 2759 0 2801
rect -270 2641 -258 2759
rect -140 2641 0 2759
rect -270 2599 0 2641
rect -270 2481 -258 2599
rect -140 2481 0 2599
rect -270 2439 0 2481
rect -270 2321 -258 2439
rect -140 2321 0 2439
rect -270 2279 0 2321
rect -270 2161 -258 2279
rect -140 2161 0 2279
rect -270 2119 0 2161
rect -270 2001 -258 2119
rect -140 2001 0 2119
rect -270 1959 0 2001
rect -270 1841 -258 1959
rect -140 1841 0 1959
rect -270 1799 0 1841
rect -270 1681 -258 1799
rect -140 1681 0 1799
rect -270 1639 0 1681
rect -270 1521 -258 1639
rect -140 1521 0 1639
rect -270 1479 0 1521
rect -270 1361 -258 1479
rect -140 1361 0 1479
rect -270 1319 0 1361
rect -270 1201 -258 1319
rect -140 1201 0 1319
rect -270 1159 0 1201
rect -270 1041 -258 1159
rect -140 1041 0 1159
rect -270 999 0 1041
rect -270 881 -258 999
rect -140 881 0 999
rect -270 839 0 881
rect -270 721 -258 839
rect -140 721 0 839
rect -270 679 0 721
rect -270 561 -258 679
rect -140 561 0 679
rect -270 519 0 561
rect -270 401 -258 519
rect -140 401 0 519
rect -270 359 0 401
rect -270 241 -258 359
rect -140 241 0 359
rect -270 199 0 241
rect -270 81 -258 199
rect -140 81 0 199
rect -270 39 0 81
rect -270 -79 -258 39
rect -140 0 0 39
rect 6000 6961 6140 7000
rect 6258 6961 6270 7079
rect 6000 6919 6270 6961
rect 6000 6801 6140 6919
rect 6258 6801 6270 6919
rect 6000 6759 6270 6801
rect 6000 6641 6140 6759
rect 6258 6641 6270 6759
rect 6000 6599 6270 6641
rect 6000 6481 6140 6599
rect 6258 6481 6270 6599
rect 6000 6439 6270 6481
rect 6000 6321 6140 6439
rect 6258 6321 6270 6439
rect 6000 6279 6270 6321
rect 6000 6161 6140 6279
rect 6258 6161 6270 6279
rect 6000 6119 6270 6161
rect 6000 6001 6140 6119
rect 6258 6001 6270 6119
rect 6000 5959 6270 6001
rect 6000 5841 6140 5959
rect 6258 5841 6270 5959
rect 6000 5799 6270 5841
rect 6000 5681 6140 5799
rect 6258 5681 6270 5799
rect 6000 5639 6270 5681
rect 6000 5521 6140 5639
rect 6258 5521 6270 5639
rect 6000 5479 6270 5521
rect 6000 5361 6140 5479
rect 6258 5361 6270 5479
rect 6000 5319 6270 5361
rect 6000 5201 6140 5319
rect 6258 5201 6270 5319
rect 6000 5159 6270 5201
rect 6000 5041 6140 5159
rect 6258 5041 6270 5159
rect 6000 4999 6270 5041
rect 6000 4881 6140 4999
rect 6258 4881 6270 4999
rect 6000 4839 6270 4881
rect 6000 4721 6140 4839
rect 6258 4721 6270 4839
rect 6000 4679 6270 4721
rect 6000 4561 6140 4679
rect 6258 4561 6270 4679
rect 6000 4519 6270 4561
rect 6000 4401 6140 4519
rect 6258 4401 6270 4519
rect 6000 4359 6270 4401
rect 6000 4241 6140 4359
rect 6258 4241 6270 4359
rect 6000 4199 6270 4241
rect 6000 4081 6140 4199
rect 6258 4081 6270 4199
rect 6000 4039 6270 4081
rect 6000 3921 6140 4039
rect 6258 3921 6270 4039
rect 6000 3879 6270 3921
rect 6000 3761 6140 3879
rect 6258 3761 6270 3879
rect 6000 3719 6270 3761
rect 6000 3601 6140 3719
rect 6258 3601 6270 3719
rect 6000 3559 6270 3601
rect 6000 3441 6140 3559
rect 6258 3441 6270 3559
rect 6000 3399 6270 3441
rect 6000 3281 6140 3399
rect 6258 3281 6270 3399
rect 6000 3239 6270 3281
rect 6000 3121 6140 3239
rect 6258 3121 6270 3239
rect 6000 3079 6270 3121
rect 6000 2961 6140 3079
rect 6258 2961 6270 3079
rect 6000 2919 6270 2961
rect 6000 2801 6140 2919
rect 6258 2801 6270 2919
rect 6000 2759 6270 2801
rect 6000 2641 6140 2759
rect 6258 2641 6270 2759
rect 6000 2599 6270 2641
rect 6000 2481 6140 2599
rect 6258 2481 6270 2599
rect 6000 2439 6270 2481
rect 6000 2321 6140 2439
rect 6258 2321 6270 2439
rect 6000 2279 6270 2321
rect 6000 2161 6140 2279
rect 6258 2161 6270 2279
rect 6000 2119 6270 2161
rect 6000 2001 6140 2119
rect 6258 2001 6270 2119
rect 6000 1959 6270 2001
rect 6000 1841 6140 1959
rect 6258 1841 6270 1959
rect 6000 1799 6270 1841
rect 6000 1681 6140 1799
rect 6258 1681 6270 1799
rect 6000 1639 6270 1681
rect 6000 1521 6140 1639
rect 6258 1521 6270 1639
rect 6000 1479 6270 1521
rect 6000 1361 6140 1479
rect 6258 1361 6270 1479
rect 6000 1319 6270 1361
rect 6000 1201 6140 1319
rect 6258 1201 6270 1319
rect 6000 1159 6270 1201
rect 6000 1041 6140 1159
rect 6258 1041 6270 1159
rect 6000 999 6270 1041
rect 6000 881 6140 999
rect 6258 881 6270 999
rect 6000 839 6270 881
rect 6000 721 6140 839
rect 6258 721 6270 839
rect 6000 679 6270 721
rect 6000 561 6140 679
rect 6258 561 6270 679
rect 6000 519 6270 561
rect 6000 401 6140 519
rect 6258 401 6270 519
rect 6000 359 6270 401
rect 6000 241 6140 359
rect 6258 241 6270 359
rect 6000 199 6270 241
rect 6000 81 6140 199
rect 6258 81 6270 199
rect 6000 39 6270 81
rect 6000 0 6140 39
rect -140 -79 6140 0
rect 6258 -79 6270 39
rect -270 -140 6270 -79
rect -270 -258 -258 -140
rect -140 -258 -19 -140
rect 99 -258 141 -140
rect 259 -258 301 -140
rect 419 -258 461 -140
rect 579 -258 621 -140
rect 739 -258 781 -140
rect 899 -258 941 -140
rect 1059 -258 1101 -140
rect 1219 -258 1261 -140
rect 1379 -258 1421 -140
rect 1539 -258 1581 -140
rect 1699 -258 1741 -140
rect 1859 -258 1901 -140
rect 2019 -258 2061 -140
rect 2179 -258 2221 -140
rect 2339 -258 2381 -140
rect 2499 -258 2541 -140
rect 2659 -258 2701 -140
rect 2819 -258 2861 -140
rect 2979 -258 3021 -140
rect 3139 -258 3181 -140
rect 3299 -258 3341 -140
rect 3459 -258 3501 -140
rect 3619 -258 3661 -140
rect 3779 -258 3821 -140
rect 3939 -258 3981 -140
rect 4099 -258 4141 -140
rect 4259 -258 4301 -140
rect 4419 -258 4461 -140
rect 4579 -258 4621 -140
rect 4739 -258 4781 -140
rect 4899 -258 4941 -140
rect 5059 -258 5101 -140
rect 5219 -258 5261 -140
rect 5379 -258 5421 -140
rect 5539 -258 5581 -140
rect 5699 -258 5741 -140
rect 5859 -258 5901 -140
rect 6019 -258 6140 -140
rect 6258 -258 6270 -140
rect -270 -270 6270 -258
<< via4 >>
rect -258 7140 -140 7258
rect -19 7140 99 7258
rect 141 7140 259 7258
rect 301 7140 419 7258
rect 461 7140 579 7258
rect 621 7140 739 7258
rect 781 7140 899 7258
rect 941 7140 1059 7258
rect 1101 7140 1219 7258
rect 1261 7140 1379 7258
rect 1421 7140 1539 7258
rect 1581 7140 1699 7258
rect 1741 7140 1859 7258
rect 1901 7140 2019 7258
rect 2061 7140 2179 7258
rect 2221 7140 2339 7258
rect 2381 7140 2499 7258
rect 2541 7140 2659 7258
rect 2701 7140 2819 7258
rect 2861 7140 2979 7258
rect 3021 7140 3139 7258
rect 3181 7140 3299 7258
rect 3341 7140 3459 7258
rect 3501 7140 3619 7258
rect 3661 7140 3779 7258
rect 3821 7140 3939 7258
rect 3981 7140 4099 7258
rect 4141 7140 4259 7258
rect 4301 7140 4419 7258
rect 4461 7140 4579 7258
rect 4621 7140 4739 7258
rect 4781 7140 4899 7258
rect 4941 7140 5059 7258
rect 5101 7140 5219 7258
rect 5261 7140 5379 7258
rect 5421 7140 5539 7258
rect 5581 7140 5699 7258
rect 5741 7140 5859 7258
rect 5901 7140 6019 7258
rect 6140 7140 6258 7258
rect -258 6961 -140 7079
rect -258 6801 -140 6919
rect -258 6641 -140 6759
rect -258 6481 -140 6599
rect -258 6321 -140 6439
rect -258 6161 -140 6279
rect -258 6001 -140 6119
rect -258 5841 -140 5959
rect -258 5681 -140 5799
rect -258 5521 -140 5639
rect -258 5361 -140 5479
rect -258 5201 -140 5319
rect -258 5041 -140 5159
rect -258 4881 -140 4999
rect -258 4721 -140 4839
rect -258 4561 -140 4679
rect -258 4401 -140 4519
rect -258 4241 -140 4359
rect -258 4081 -140 4199
rect -258 3921 -140 4039
rect -258 3761 -140 3879
rect -258 3601 -140 3719
rect -258 3441 -140 3559
rect -258 3281 -140 3399
rect -258 3121 -140 3239
rect -258 2961 -140 3079
rect -258 2801 -140 2919
rect -258 2641 -140 2759
rect -258 2481 -140 2599
rect -258 2321 -140 2439
rect -258 2161 -140 2279
rect -258 2001 -140 2119
rect -258 1841 -140 1959
rect -258 1681 -140 1799
rect -258 1521 -140 1639
rect -258 1361 -140 1479
rect -258 1201 -140 1319
rect -258 1041 -140 1159
rect -258 881 -140 999
rect -258 721 -140 839
rect -258 561 -140 679
rect -258 401 -140 519
rect -258 241 -140 359
rect -258 81 -140 199
rect -258 -79 -140 39
rect 6140 6961 6258 7079
rect 6140 6801 6258 6919
rect 6140 6641 6258 6759
rect 6140 6481 6258 6599
rect 6140 6321 6258 6439
rect 6140 6161 6258 6279
rect 6140 6001 6258 6119
rect 6140 5841 6258 5959
rect 6140 5681 6258 5799
rect 6140 5521 6258 5639
rect 6140 5361 6258 5479
rect 6140 5201 6258 5319
rect 6140 5041 6258 5159
rect 6140 4881 6258 4999
rect 6140 4721 6258 4839
rect 6140 4561 6258 4679
rect 6140 4401 6258 4519
rect 6140 4241 6258 4359
rect 6140 4081 6258 4199
rect 6140 3921 6258 4039
rect 6140 3761 6258 3879
rect 6140 3601 6258 3719
rect 6140 3441 6258 3559
rect 6140 3281 6258 3399
rect 6140 3121 6258 3239
rect 6140 2961 6258 3079
rect 6140 2801 6258 2919
rect 6140 2641 6258 2759
rect 6140 2481 6258 2599
rect 6140 2321 6258 2439
rect 6140 2161 6258 2279
rect 6140 2001 6258 2119
rect 6140 1841 6258 1959
rect 6140 1681 6258 1799
rect 6140 1521 6258 1639
rect 6140 1361 6258 1479
rect 6140 1201 6258 1319
rect 6140 1041 6258 1159
rect 6140 881 6258 999
rect 6140 721 6258 839
rect 6140 561 6258 679
rect 6140 401 6258 519
rect 6140 241 6258 359
rect 6140 81 6258 199
rect 6140 -79 6258 39
rect -258 -258 -140 -140
rect -19 -258 99 -140
rect 141 -258 259 -140
rect 301 -258 419 -140
rect 461 -258 579 -140
rect 621 -258 739 -140
rect 781 -258 899 -140
rect 941 -258 1059 -140
rect 1101 -258 1219 -140
rect 1261 -258 1379 -140
rect 1421 -258 1539 -140
rect 1581 -258 1699 -140
rect 1741 -258 1859 -140
rect 1901 -258 2019 -140
rect 2061 -258 2179 -140
rect 2221 -258 2339 -140
rect 2381 -258 2499 -140
rect 2541 -258 2659 -140
rect 2701 -258 2819 -140
rect 2861 -258 2979 -140
rect 3021 -258 3139 -140
rect 3181 -258 3299 -140
rect 3341 -258 3459 -140
rect 3501 -258 3619 -140
rect 3661 -258 3779 -140
rect 3821 -258 3939 -140
rect 3981 -258 4099 -140
rect 4141 -258 4259 -140
rect 4301 -258 4419 -140
rect 4461 -258 4579 -140
rect 4621 -258 4739 -140
rect 4781 -258 4899 -140
rect 4941 -258 5059 -140
rect 5101 -258 5219 -140
rect 5261 -258 5379 -140
rect 5421 -258 5539 -140
rect 5581 -258 5699 -140
rect 5741 -258 5859 -140
rect 5901 -258 6019 -140
rect 6140 -258 6258 -140
<< metal5 >>
rect -270 7258 6270 7270
rect -270 7140 -258 7258
rect -140 7140 -19 7258
rect 99 7140 141 7258
rect 259 7140 301 7258
rect 419 7140 461 7258
rect 579 7140 621 7258
rect 739 7140 781 7258
rect 899 7140 941 7258
rect 1059 7140 1101 7258
rect 1219 7140 1261 7258
rect 1379 7140 1421 7258
rect 1539 7140 1581 7258
rect 1699 7140 1741 7258
rect 1859 7140 1901 7258
rect 2019 7140 2061 7258
rect 2179 7140 2221 7258
rect 2339 7140 2381 7258
rect 2499 7140 2541 7258
rect 2659 7140 2701 7258
rect 2819 7140 2861 7258
rect 2979 7140 3021 7258
rect 3139 7140 3181 7258
rect 3299 7140 3341 7258
rect 3459 7140 3501 7258
rect 3619 7140 3661 7258
rect 3779 7140 3821 7258
rect 3939 7140 3981 7258
rect 4099 7140 4141 7258
rect 4259 7140 4301 7258
rect 4419 7140 4461 7258
rect 4579 7140 4621 7258
rect 4739 7140 4781 7258
rect 4899 7140 4941 7258
rect 5059 7140 5101 7258
rect 5219 7140 5261 7258
rect 5379 7140 5421 7258
rect 5539 7140 5581 7258
rect 5699 7140 5741 7258
rect 5859 7140 5901 7258
rect 6019 7140 6140 7258
rect 6258 7140 6270 7258
rect -270 7079 6270 7140
rect -270 6961 -258 7079
rect -140 6961 6140 7079
rect 6258 6961 6270 7079
rect -270 6919 6270 6961
rect -270 6801 -258 6919
rect -140 6801 6140 6919
rect 6258 6801 6270 6919
rect -270 6759 6270 6801
rect -270 6641 -258 6759
rect -140 6641 6140 6759
rect 6258 6641 6270 6759
rect -270 6599 6270 6641
rect -270 6481 -258 6599
rect -140 6481 6140 6599
rect 6258 6481 6270 6599
rect -270 6439 6270 6481
rect -270 6321 -258 6439
rect -140 6321 6140 6439
rect 6258 6321 6270 6439
rect -270 6279 6270 6321
rect -270 6161 -258 6279
rect -140 6161 6140 6279
rect 6258 6161 6270 6279
rect -270 6119 6270 6161
rect -270 6001 -258 6119
rect -140 6001 6140 6119
rect 6258 6001 6270 6119
rect -270 5959 6270 6001
rect -270 5841 -258 5959
rect -140 5841 6140 5959
rect 6258 5841 6270 5959
rect -270 5799 6270 5841
rect -270 5681 -258 5799
rect -140 5681 6140 5799
rect 6258 5681 6270 5799
rect -270 5639 6270 5681
rect -270 5521 -258 5639
rect -140 5521 6140 5639
rect 6258 5521 6270 5639
rect -270 5479 6270 5521
rect -270 5361 -258 5479
rect -140 5361 6140 5479
rect 6258 5361 6270 5479
rect -270 5319 6270 5361
rect -270 5201 -258 5319
rect -140 5201 6140 5319
rect 6258 5201 6270 5319
rect -270 5159 6270 5201
rect -270 5041 -258 5159
rect -140 5041 6140 5159
rect 6258 5041 6270 5159
rect -270 4999 6270 5041
rect -270 4881 -258 4999
rect -140 4881 6140 4999
rect 6258 4881 6270 4999
rect -270 4839 6270 4881
rect -270 4721 -258 4839
rect -140 4721 6140 4839
rect 6258 4721 6270 4839
rect -270 4679 6270 4721
rect -270 4561 -258 4679
rect -140 4561 6140 4679
rect 6258 4561 6270 4679
rect -270 4519 6270 4561
rect -270 4401 -258 4519
rect -140 4401 6140 4519
rect 6258 4401 6270 4519
rect -270 4359 6270 4401
rect -270 4241 -258 4359
rect -140 4241 6140 4359
rect 6258 4241 6270 4359
rect -270 4199 6270 4241
rect -270 4081 -258 4199
rect -140 4081 6140 4199
rect 6258 4081 6270 4199
rect -270 4039 6270 4081
rect -270 3921 -258 4039
rect -140 3921 6140 4039
rect 6258 3921 6270 4039
rect -270 3879 6270 3921
rect -270 3761 -258 3879
rect -140 3761 6140 3879
rect 6258 3761 6270 3879
rect -270 3719 6270 3761
rect -270 3601 -258 3719
rect -140 3601 6140 3719
rect 6258 3601 6270 3719
rect -270 3559 6270 3601
rect -270 3441 -258 3559
rect -140 3441 6140 3559
rect 6258 3441 6270 3559
rect -270 3399 6270 3441
rect -270 3281 -258 3399
rect -140 3281 6140 3399
rect 6258 3281 6270 3399
rect -270 3239 6270 3281
rect -270 3121 -258 3239
rect -140 3121 6140 3239
rect 6258 3121 6270 3239
rect -270 3079 6270 3121
rect -270 2961 -258 3079
rect -140 2961 6140 3079
rect 6258 2961 6270 3079
rect -270 2919 6270 2961
rect -270 2801 -258 2919
rect -140 2801 6140 2919
rect 6258 2801 6270 2919
rect -270 2759 6270 2801
rect -270 2641 -258 2759
rect -140 2641 6140 2759
rect 6258 2641 6270 2759
rect -270 2599 6270 2641
rect -270 2481 -258 2599
rect -140 2481 6140 2599
rect 6258 2481 6270 2599
rect -270 2439 6270 2481
rect -270 2321 -258 2439
rect -140 2321 6140 2439
rect 6258 2321 6270 2439
rect -270 2279 6270 2321
rect -270 2161 -258 2279
rect -140 2161 6140 2279
rect 6258 2161 6270 2279
rect -270 2119 6270 2161
rect -270 2001 -258 2119
rect -140 2001 6140 2119
rect 6258 2001 6270 2119
rect -270 1959 6270 2001
rect -270 1841 -258 1959
rect -140 1841 6140 1959
rect 6258 1841 6270 1959
rect -270 1799 6270 1841
rect -270 1681 -258 1799
rect -140 1681 6140 1799
rect 6258 1681 6270 1799
rect -270 1639 6270 1681
rect -270 1521 -258 1639
rect -140 1521 6140 1639
rect 6258 1521 6270 1639
rect -270 1479 6270 1521
rect -270 1361 -258 1479
rect -140 1361 6140 1479
rect 6258 1361 6270 1479
rect -270 1319 6270 1361
rect -270 1201 -258 1319
rect -140 1201 6140 1319
rect 6258 1201 6270 1319
rect -270 1159 6270 1201
rect -270 1041 -258 1159
rect -140 1041 6140 1159
rect 6258 1041 6270 1159
rect -270 999 6270 1041
rect -270 881 -258 999
rect -140 881 6140 999
rect 6258 881 6270 999
rect -270 839 6270 881
rect -270 721 -258 839
rect -140 721 6140 839
rect 6258 721 6270 839
rect -270 679 6270 721
rect -270 561 -258 679
rect -140 561 6140 679
rect 6258 561 6270 679
rect -270 519 6270 561
rect -270 401 -258 519
rect -140 401 6140 519
rect 6258 401 6270 519
rect -270 359 6270 401
rect -270 241 -258 359
rect -140 241 6140 359
rect 6258 241 6270 359
rect -270 199 6270 241
rect -270 81 -258 199
rect -140 81 6140 199
rect 6258 81 6270 199
rect -270 39 6270 81
rect -270 -79 -258 39
rect -140 -79 6140 39
rect 6258 -79 6270 39
rect -270 -140 6270 -79
rect -270 -258 -258 -140
rect -140 -258 -19 -140
rect 99 -258 141 -140
rect 259 -258 301 -140
rect 419 -258 461 -140
rect 579 -258 621 -140
rect 739 -258 781 -140
rect 899 -258 941 -140
rect 1059 -258 1101 -140
rect 1219 -258 1261 -140
rect 1379 -258 1421 -140
rect 1539 -258 1581 -140
rect 1699 -258 1741 -140
rect 1859 -258 1901 -140
rect 2019 -258 2061 -140
rect 2179 -258 2221 -140
rect 2339 -258 2381 -140
rect 2499 -258 2541 -140
rect 2659 -258 2701 -140
rect 2819 -258 2861 -140
rect 2979 -258 3021 -140
rect 3139 -258 3181 -140
rect 3299 -258 3341 -140
rect 3459 -258 3501 -140
rect 3619 -258 3661 -140
rect 3779 -258 3821 -140
rect 3939 -258 3981 -140
rect 4099 -258 4141 -140
rect 4259 -258 4301 -140
rect 4419 -258 4461 -140
rect 4579 -258 4621 -140
rect 4739 -258 4781 -140
rect 4899 -258 4941 -140
rect 5059 -258 5101 -140
rect 5219 -258 5261 -140
rect 5379 -258 5421 -140
rect 5539 -258 5581 -140
rect 5699 -258 5741 -140
rect 5859 -258 5901 -140
rect 6019 -258 6140 -140
rect 6258 -258 6270 -140
rect -270 -270 6270 -258
<< glass >>
rect 0 0 6000 7000
<< labels >>
flabel metal5 s -140 -140 6140 7140 0 FreeSans 1000 0 0 0 PAD
port 1 nsew
<< properties >>
string GDS_END 11530
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_ef_io__bare_pad.gds
string GDS_START 134
<< end >>
