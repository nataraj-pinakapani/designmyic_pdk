magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 8 5 8 9 6 C0
port 1 nsew
rlabel  s 8 0 8 4 6 C0
port 1 nsew
rlabel  s 7 7 7 9 6 C0
port 1 nsew
rlabel  s 7 5 7 6 6 C0
port 1 nsew
rlabel  s 7 3 7 4 6 C0
port 1 nsew
rlabel  s 7 0 7 2 6 C0
port 1 nsew
rlabel  s 5 7 6 9 6 C0
port 1 nsew
rlabel  s 5 5 6 6 6 C0
port 1 nsew
rlabel  s 5 3 6 4 6 C0
port 1 nsew
rlabel  s 5 0 6 2 6 C0
port 1 nsew
rlabel  s 4 5 4 9 6 C0
port 1 nsew
rlabel  s 4 0 4 4 6 C0
port 1 nsew
rlabel  s 3 7 3 9 6 C0
port 1 nsew
rlabel  s 3 5 3 6 6 C0
port 1 nsew
rlabel  s 3 3 3 4 6 C0
port 1 nsew
rlabel  s 3 0 3 2 6 C0
port 1 nsew
rlabel  s 1 7 2 9 6 C0
port 1 nsew
rlabel  s 1 5 2 6 6 C0
port 1 nsew
rlabel  s 1 3 2 4 6 C0
port 1 nsew
rlabel  s 1 0 2 2 6 C0
port 1 nsew
rlabel  s 0 9 8 9 6 C0
port 1 nsew
rlabel  s 0 5 0 9 4 C0
port 1 nsew
rlabel  s 0 4 8 5 6 C0
port 1 nsew
rlabel  s 0 0 0 4 4 C0
port 1 nsew
rlabel  s 0 0 8 0 8 C0
port 1 nsew
rlabel  s 8 7 8 8 6 C1
port 2 nsew
rlabel  s 8 5 8 6 6 C1
port 2 nsew
rlabel  s 8 2 8 4 6 C1
port 2 nsew
rlabel  s 8 1 8 2 6 C1
port 2 nsew
rlabel  s 6 7 6 8 6 C1
port 2 nsew
rlabel  s 6 5 6 6 6 C1
port 2 nsew
rlabel  s 6 2 6 4 6 C1
port 2 nsew
rlabel  s 6 1 6 2 6 C1
port 2 nsew
rlabel  s 5 7 5 8 6 C1
port 2 nsew
rlabel  s 5 6 8 7 6 C1
port 2 nsew
rlabel  s 5 5 5 6 6 C1
port 2 nsew
rlabel  s 5 2 5 4 6 C1
port 2 nsew
rlabel  s 5 2 8 2 6 C1
port 2 nsew
rlabel  s 5 1 5 2 6 C1
port 2 nsew
rlabel  s 3 7 4 8 6 C1
port 2 nsew
rlabel  s 3 5 4 6 6 C1
port 2 nsew
rlabel  s 3 2 4 4 6 C1
port 2 nsew
rlabel  s 3 1 4 2 6 C1
port 2 nsew
rlabel  s 2 7 2 8 6 C1
port 2 nsew
rlabel  s 2 5 2 6 6 C1
port 2 nsew
rlabel  s 2 2 2 4 6 C1
port 2 nsew
rlabel  s 2 1 2 2 6 C1
port 2 nsew
rlabel  s 1 7 1 8 6 C1
port 2 nsew
rlabel  s 1 6 4 7 6 C1
port 2 nsew
rlabel  s 1 5 1 6 6 C1
port 2 nsew
rlabel  s 1 2 1 4 6 C1
port 2 nsew
rlabel  s 1 2 4 2 6 C1
port 2 nsew
rlabel  s 1 1 1 2 6 C1
port 2 nsew
rlabel r s 0 0 8 9 6 M5
port 3 nsew
rlabel metal_blue s 6 6 6 6 6 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 8 9
string LEFview TRUE
<< end >>
