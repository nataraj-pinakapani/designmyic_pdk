magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 258 -30 3550 992
<< pwell >>
rect -36 1052 3501 1138
rect -36 -90 50 1052
rect -36 -176 3493 -90
<< mvpmos >>
rect 756 665 1756 765
rect 1886 665 3286 765
rect 756 509 1756 609
rect 1886 509 3286 609
rect 756 353 1756 453
rect 1886 353 3286 453
rect 756 197 1756 297
rect 1886 197 3286 297
<< mvpdiff >>
rect 756 810 1756 818
rect 756 776 826 810
rect 860 776 894 810
rect 928 776 962 810
rect 996 776 1030 810
rect 1064 776 1098 810
rect 1132 776 1166 810
rect 1200 776 1234 810
rect 1268 776 1302 810
rect 1336 776 1370 810
rect 1404 776 1438 810
rect 1472 776 1506 810
rect 1540 776 1574 810
rect 1608 776 1642 810
rect 1676 776 1710 810
rect 1744 776 1756 810
rect 756 765 1756 776
rect 1886 810 3286 818
rect 1886 776 1948 810
rect 1982 776 2016 810
rect 2050 776 2084 810
rect 2118 776 2152 810
rect 2186 776 2220 810
rect 2254 776 2288 810
rect 2322 776 2356 810
rect 2390 776 2424 810
rect 2458 776 2492 810
rect 2526 776 2560 810
rect 2594 776 2628 810
rect 2662 776 2696 810
rect 2730 776 2764 810
rect 2798 776 2832 810
rect 2866 776 2900 810
rect 2934 776 2968 810
rect 3002 776 3036 810
rect 3070 776 3104 810
rect 3138 776 3172 810
rect 3206 776 3240 810
rect 3274 776 3286 810
rect 1886 765 3286 776
rect 756 654 1756 665
rect 756 620 826 654
rect 860 620 894 654
rect 928 620 962 654
rect 996 620 1030 654
rect 1064 620 1098 654
rect 1132 620 1166 654
rect 1200 620 1234 654
rect 1268 620 1302 654
rect 1336 620 1370 654
rect 1404 620 1438 654
rect 1472 620 1506 654
rect 1540 620 1574 654
rect 1608 620 1642 654
rect 1676 620 1710 654
rect 1744 620 1756 654
rect 756 609 1756 620
rect 1886 654 3286 665
rect 1886 620 1948 654
rect 1982 620 2016 654
rect 2050 620 2084 654
rect 2118 620 2152 654
rect 2186 620 2220 654
rect 2254 620 2288 654
rect 2322 620 2356 654
rect 2390 620 2424 654
rect 2458 620 2492 654
rect 2526 620 2560 654
rect 2594 620 2628 654
rect 2662 620 2696 654
rect 2730 620 2764 654
rect 2798 620 2832 654
rect 2866 620 2900 654
rect 2934 620 2968 654
rect 3002 620 3036 654
rect 3070 620 3104 654
rect 3138 620 3172 654
rect 3206 620 3240 654
rect 3274 620 3286 654
rect 1886 609 3286 620
rect 756 498 1756 509
rect 756 464 826 498
rect 860 464 894 498
rect 928 464 962 498
rect 996 464 1030 498
rect 1064 464 1098 498
rect 1132 464 1166 498
rect 1200 464 1234 498
rect 1268 464 1302 498
rect 1336 464 1370 498
rect 1404 464 1438 498
rect 1472 464 1506 498
rect 1540 464 1574 498
rect 1608 464 1642 498
rect 1676 464 1710 498
rect 1744 464 1756 498
rect 756 453 1756 464
rect 1886 498 3286 509
rect 1886 464 1948 498
rect 1982 464 2016 498
rect 2050 464 2084 498
rect 2118 464 2152 498
rect 2186 464 2220 498
rect 2254 464 2288 498
rect 2322 464 2356 498
rect 2390 464 2424 498
rect 2458 464 2492 498
rect 2526 464 2560 498
rect 2594 464 2628 498
rect 2662 464 2696 498
rect 2730 464 2764 498
rect 2798 464 2832 498
rect 2866 464 2900 498
rect 2934 464 2968 498
rect 3002 464 3036 498
rect 3070 464 3104 498
rect 3138 464 3172 498
rect 3206 464 3240 498
rect 3274 464 3286 498
rect 1886 453 3286 464
rect 756 342 1756 353
rect 756 308 826 342
rect 860 308 894 342
rect 928 308 962 342
rect 996 308 1030 342
rect 1064 308 1098 342
rect 1132 308 1166 342
rect 1200 308 1234 342
rect 1268 308 1302 342
rect 1336 308 1370 342
rect 1404 308 1438 342
rect 1472 308 1506 342
rect 1540 308 1574 342
rect 1608 308 1642 342
rect 1676 308 1710 342
rect 1744 308 1756 342
rect 756 297 1756 308
rect 1886 342 3286 353
rect 1886 308 1948 342
rect 1982 308 2016 342
rect 2050 308 2084 342
rect 2118 308 2152 342
rect 2186 308 2220 342
rect 2254 308 2288 342
rect 2322 308 2356 342
rect 2390 308 2424 342
rect 2458 308 2492 342
rect 2526 308 2560 342
rect 2594 308 2628 342
rect 2662 308 2696 342
rect 2730 308 2764 342
rect 2798 308 2832 342
rect 2866 308 2900 342
rect 2934 308 2968 342
rect 3002 308 3036 342
rect 3070 308 3104 342
rect 3138 308 3172 342
rect 3206 308 3240 342
rect 3274 308 3286 342
rect 1886 297 3286 308
rect 756 186 1756 197
rect 756 152 826 186
rect 860 152 894 186
rect 928 152 962 186
rect 996 152 1030 186
rect 1064 152 1098 186
rect 1132 152 1166 186
rect 1200 152 1234 186
rect 1268 152 1302 186
rect 1336 152 1370 186
rect 1404 152 1438 186
rect 1472 152 1506 186
rect 1540 152 1574 186
rect 1608 152 1642 186
rect 1676 152 1710 186
rect 1744 152 1756 186
rect 756 144 1756 152
rect 1886 186 3286 197
rect 1886 152 1948 186
rect 1982 152 2016 186
rect 2050 152 2084 186
rect 2118 152 2152 186
rect 2186 152 2220 186
rect 2254 152 2288 186
rect 2322 152 2356 186
rect 2390 152 2424 186
rect 2458 152 2492 186
rect 2526 152 2560 186
rect 2594 152 2628 186
rect 2662 152 2696 186
rect 2730 152 2764 186
rect 2798 152 2832 186
rect 2866 152 2900 186
rect 2934 152 2968 186
rect 3002 152 3036 186
rect 3070 152 3104 186
rect 3138 152 3172 186
rect 3206 152 3240 186
rect 3274 152 3286 186
rect 1886 144 3286 152
<< mvpdiffc >>
rect 826 776 860 810
rect 894 776 928 810
rect 962 776 996 810
rect 1030 776 1064 810
rect 1098 776 1132 810
rect 1166 776 1200 810
rect 1234 776 1268 810
rect 1302 776 1336 810
rect 1370 776 1404 810
rect 1438 776 1472 810
rect 1506 776 1540 810
rect 1574 776 1608 810
rect 1642 776 1676 810
rect 1710 776 1744 810
rect 1948 776 1982 810
rect 2016 776 2050 810
rect 2084 776 2118 810
rect 2152 776 2186 810
rect 2220 776 2254 810
rect 2288 776 2322 810
rect 2356 776 2390 810
rect 2424 776 2458 810
rect 2492 776 2526 810
rect 2560 776 2594 810
rect 2628 776 2662 810
rect 2696 776 2730 810
rect 2764 776 2798 810
rect 2832 776 2866 810
rect 2900 776 2934 810
rect 2968 776 3002 810
rect 3036 776 3070 810
rect 3104 776 3138 810
rect 3172 776 3206 810
rect 3240 776 3274 810
rect 826 620 860 654
rect 894 620 928 654
rect 962 620 996 654
rect 1030 620 1064 654
rect 1098 620 1132 654
rect 1166 620 1200 654
rect 1234 620 1268 654
rect 1302 620 1336 654
rect 1370 620 1404 654
rect 1438 620 1472 654
rect 1506 620 1540 654
rect 1574 620 1608 654
rect 1642 620 1676 654
rect 1710 620 1744 654
rect 1948 620 1982 654
rect 2016 620 2050 654
rect 2084 620 2118 654
rect 2152 620 2186 654
rect 2220 620 2254 654
rect 2288 620 2322 654
rect 2356 620 2390 654
rect 2424 620 2458 654
rect 2492 620 2526 654
rect 2560 620 2594 654
rect 2628 620 2662 654
rect 2696 620 2730 654
rect 2764 620 2798 654
rect 2832 620 2866 654
rect 2900 620 2934 654
rect 2968 620 3002 654
rect 3036 620 3070 654
rect 3104 620 3138 654
rect 3172 620 3206 654
rect 3240 620 3274 654
rect 826 464 860 498
rect 894 464 928 498
rect 962 464 996 498
rect 1030 464 1064 498
rect 1098 464 1132 498
rect 1166 464 1200 498
rect 1234 464 1268 498
rect 1302 464 1336 498
rect 1370 464 1404 498
rect 1438 464 1472 498
rect 1506 464 1540 498
rect 1574 464 1608 498
rect 1642 464 1676 498
rect 1710 464 1744 498
rect 1948 464 1982 498
rect 2016 464 2050 498
rect 2084 464 2118 498
rect 2152 464 2186 498
rect 2220 464 2254 498
rect 2288 464 2322 498
rect 2356 464 2390 498
rect 2424 464 2458 498
rect 2492 464 2526 498
rect 2560 464 2594 498
rect 2628 464 2662 498
rect 2696 464 2730 498
rect 2764 464 2798 498
rect 2832 464 2866 498
rect 2900 464 2934 498
rect 2968 464 3002 498
rect 3036 464 3070 498
rect 3104 464 3138 498
rect 3172 464 3206 498
rect 3240 464 3274 498
rect 826 308 860 342
rect 894 308 928 342
rect 962 308 996 342
rect 1030 308 1064 342
rect 1098 308 1132 342
rect 1166 308 1200 342
rect 1234 308 1268 342
rect 1302 308 1336 342
rect 1370 308 1404 342
rect 1438 308 1472 342
rect 1506 308 1540 342
rect 1574 308 1608 342
rect 1642 308 1676 342
rect 1710 308 1744 342
rect 1948 308 1982 342
rect 2016 308 2050 342
rect 2084 308 2118 342
rect 2152 308 2186 342
rect 2220 308 2254 342
rect 2288 308 2322 342
rect 2356 308 2390 342
rect 2424 308 2458 342
rect 2492 308 2526 342
rect 2560 308 2594 342
rect 2628 308 2662 342
rect 2696 308 2730 342
rect 2764 308 2798 342
rect 2832 308 2866 342
rect 2900 308 2934 342
rect 2968 308 3002 342
rect 3036 308 3070 342
rect 3104 308 3138 342
rect 3172 308 3206 342
rect 3240 308 3274 342
rect 826 152 860 186
rect 894 152 928 186
rect 962 152 996 186
rect 1030 152 1064 186
rect 1098 152 1132 186
rect 1166 152 1200 186
rect 1234 152 1268 186
rect 1302 152 1336 186
rect 1370 152 1404 186
rect 1438 152 1472 186
rect 1506 152 1540 186
rect 1574 152 1608 186
rect 1642 152 1676 186
rect 1710 152 1744 186
rect 1948 152 1982 186
rect 2016 152 2050 186
rect 2084 152 2118 186
rect 2152 152 2186 186
rect 2220 152 2254 186
rect 2288 152 2322 186
rect 2356 152 2390 186
rect 2424 152 2458 186
rect 2492 152 2526 186
rect 2560 152 2594 186
rect 2628 152 2662 186
rect 2696 152 2730 186
rect 2764 152 2798 186
rect 2832 152 2866 186
rect 2900 152 2934 186
rect 2968 152 3002 186
rect 3036 152 3070 186
rect 3104 152 3138 186
rect 3172 152 3206 186
rect 3240 152 3274 186
<< mvpsubdiff >>
rect -10 1088 69 1112
rect 24 1078 69 1088
rect 103 1078 137 1112
rect 171 1078 205 1112
rect 239 1078 273 1112
rect 307 1078 341 1112
rect 375 1078 409 1112
rect 443 1078 477 1112
rect 511 1078 545 1112
rect 579 1078 613 1112
rect 647 1078 681 1112
rect 715 1078 749 1112
rect 783 1078 817 1112
rect 851 1078 885 1112
rect 919 1078 953 1112
rect 987 1078 1021 1112
rect 1055 1078 1089 1112
rect 1123 1078 1157 1112
rect 1191 1078 1225 1112
rect 1259 1078 1293 1112
rect 1327 1078 1361 1112
rect 1395 1078 1429 1112
rect 1463 1078 1497 1112
rect 1531 1078 1565 1112
rect 1599 1078 1633 1112
rect 1667 1078 1701 1112
rect 1735 1078 1769 1112
rect 1803 1078 1837 1112
rect 1871 1078 1905 1112
rect 1939 1078 1973 1112
rect 2007 1078 2041 1112
rect 2075 1078 2109 1112
rect 2143 1078 2177 1112
rect 2211 1078 2245 1112
rect 2279 1078 2313 1112
rect 2347 1078 2381 1112
rect 2415 1078 2449 1112
rect 2483 1078 2517 1112
rect 2551 1078 2585 1112
rect 2619 1078 2653 1112
rect 2687 1078 2721 1112
rect 2755 1078 2789 1112
rect 2823 1078 2857 1112
rect 2891 1078 2925 1112
rect 2959 1078 2993 1112
rect 3027 1078 3061 1112
rect 3095 1078 3129 1112
rect 3163 1078 3197 1112
rect 3231 1078 3265 1112
rect 3299 1078 3333 1112
rect 3367 1078 3401 1112
rect 3435 1078 3475 1112
rect -10 1020 24 1054
rect -10 952 24 986
rect -10 884 24 918
rect -10 816 24 850
rect -10 748 24 782
rect -10 680 24 714
rect -10 612 24 646
rect -10 544 24 578
rect -10 476 24 510
rect -10 408 24 442
rect -10 340 24 374
rect -10 272 24 306
rect -10 204 24 238
rect -10 136 24 170
rect -10 68 24 102
rect -10 0 24 34
rect -10 -116 24 -34
rect -10 -150 123 -116
rect 157 -150 191 -116
rect 225 -150 259 -116
rect 293 -150 327 -116
rect 361 -150 395 -116
rect 429 -150 463 -116
rect 497 -150 531 -116
rect 565 -150 599 -116
rect 633 -150 667 -116
rect 701 -150 735 -116
rect 769 -150 803 -116
rect 837 -150 871 -116
rect 905 -150 939 -116
rect 973 -150 1007 -116
rect 1041 -150 1075 -116
rect 1109 -150 3467 -116
<< mvnsubdiff >>
rect 324 892 348 926
rect 382 892 416 926
rect 450 892 484 926
rect 518 892 655 926
rect 689 892 723 926
rect 757 892 791 926
rect 825 892 859 926
rect 893 892 927 926
rect 961 892 995 926
rect 1029 892 1063 926
rect 1097 892 1131 926
rect 1165 892 1199 926
rect 1233 892 1267 926
rect 1301 892 1335 926
rect 1369 892 1403 926
rect 1437 892 1471 926
rect 1505 892 1539 926
rect 1573 892 1607 926
rect 1641 892 1675 926
rect 1709 892 1743 926
rect 1777 892 1811 926
rect 1845 892 1879 926
rect 1913 892 1947 926
rect 1981 892 2015 926
rect 2049 892 2083 926
rect 2117 892 2151 926
rect 2185 892 2219 926
rect 2253 892 2287 926
rect 2321 892 2355 926
rect 2389 892 2423 926
rect 2457 892 2491 926
rect 2525 892 2559 926
rect 2593 892 2627 926
rect 2661 892 2695 926
rect 2729 892 2763 926
rect 2797 892 2831 926
rect 2865 892 2899 926
rect 2933 892 2967 926
rect 3001 892 3035 926
rect 3069 892 3103 926
rect 3137 892 3171 926
rect 3205 892 3239 926
rect 3273 892 3307 926
rect 3341 892 3375 926
rect 3409 902 3484 926
rect 3409 892 3450 902
rect 324 842 575 892
rect 358 824 575 842
rect 358 808 393 824
rect 324 790 393 808
rect 427 790 467 824
rect 501 790 541 824
rect 3450 834 3484 868
rect 324 774 575 790
rect 358 751 575 774
rect 3450 766 3484 800
rect 358 740 393 751
rect 324 717 393 740
rect 427 717 467 751
rect 501 717 541 751
rect 324 706 575 717
rect 358 678 575 706
rect 358 672 393 678
rect 324 644 393 672
rect 427 644 467 678
rect 501 644 541 678
rect 324 638 575 644
rect 358 605 575 638
rect 358 604 393 605
rect 324 571 393 604
rect 427 571 467 605
rect 501 571 541 605
rect 324 570 575 571
rect 358 536 575 570
rect 324 532 575 536
rect 324 502 393 532
rect 358 498 393 502
rect 427 498 467 532
rect 501 498 541 532
rect 358 468 575 498
rect 324 459 575 468
rect 324 434 393 459
rect 358 425 393 434
rect 427 425 467 459
rect 501 425 541 459
rect 358 400 575 425
rect 324 386 575 400
rect 324 366 393 386
rect 358 352 393 366
rect 427 352 467 386
rect 501 352 541 386
rect 358 332 575 352
rect 324 312 575 332
rect 324 298 393 312
rect 358 278 393 298
rect 427 278 467 312
rect 501 278 541 312
rect 358 264 575 278
rect 324 238 575 264
rect 324 230 393 238
rect 358 204 393 230
rect 427 204 467 238
rect 501 204 541 238
rect 358 196 575 204
rect 3450 698 3484 732
rect 3450 630 3484 664
rect 3450 562 3484 596
rect 3450 494 3484 528
rect 3450 426 3484 460
rect 3450 358 3484 392
rect 3450 290 3484 324
rect 3450 222 3484 256
rect 324 164 575 196
rect 324 162 393 164
rect 358 130 393 162
rect 427 130 467 164
rect 501 130 541 164
rect 3450 154 3484 188
rect 358 128 575 130
rect 324 94 575 128
rect 358 70 575 94
rect 3450 70 3484 120
rect 358 60 434 70
rect 324 36 434 60
rect 468 36 502 70
rect 536 36 570 70
rect 604 36 638 70
rect 672 36 706 70
rect 740 36 774 70
rect 808 36 842 70
rect 876 36 910 70
rect 944 36 978 70
rect 1012 36 1046 70
rect 1080 36 1114 70
rect 1148 36 1182 70
rect 1216 36 1250 70
rect 1284 36 1318 70
rect 1352 36 1386 70
rect 1420 36 1454 70
rect 1488 36 1522 70
rect 1556 36 1590 70
rect 1624 36 1658 70
rect 1692 36 1726 70
rect 1760 36 1794 70
rect 1828 36 1862 70
rect 1896 36 1930 70
rect 1964 36 1998 70
rect 2032 36 2066 70
rect 2100 36 2134 70
rect 2168 36 2202 70
rect 2236 36 2270 70
rect 2304 36 2338 70
rect 2372 36 2406 70
rect 2440 36 2474 70
rect 2508 36 2542 70
rect 2576 36 2610 70
rect 2644 36 2678 70
rect 2712 36 2746 70
rect 2780 36 2814 70
rect 2848 36 2882 70
rect 2916 36 2950 70
rect 2984 36 3018 70
rect 3052 36 3086 70
rect 3120 36 3154 70
rect 3188 36 3222 70
rect 3256 36 3290 70
rect 3324 36 3358 70
rect 3392 36 3426 70
rect 3460 36 3484 70
<< mvpsubdiffcont >>
rect -10 1054 24 1088
rect 69 1078 103 1112
rect 137 1078 171 1112
rect 205 1078 239 1112
rect 273 1078 307 1112
rect 341 1078 375 1112
rect 409 1078 443 1112
rect 477 1078 511 1112
rect 545 1078 579 1112
rect 613 1078 647 1112
rect 681 1078 715 1112
rect 749 1078 783 1112
rect 817 1078 851 1112
rect 885 1078 919 1112
rect 953 1078 987 1112
rect 1021 1078 1055 1112
rect 1089 1078 1123 1112
rect 1157 1078 1191 1112
rect 1225 1078 1259 1112
rect 1293 1078 1327 1112
rect 1361 1078 1395 1112
rect 1429 1078 1463 1112
rect 1497 1078 1531 1112
rect 1565 1078 1599 1112
rect 1633 1078 1667 1112
rect 1701 1078 1735 1112
rect 1769 1078 1803 1112
rect 1837 1078 1871 1112
rect 1905 1078 1939 1112
rect 1973 1078 2007 1112
rect 2041 1078 2075 1112
rect 2109 1078 2143 1112
rect 2177 1078 2211 1112
rect 2245 1078 2279 1112
rect 2313 1078 2347 1112
rect 2381 1078 2415 1112
rect 2449 1078 2483 1112
rect 2517 1078 2551 1112
rect 2585 1078 2619 1112
rect 2653 1078 2687 1112
rect 2721 1078 2755 1112
rect 2789 1078 2823 1112
rect 2857 1078 2891 1112
rect 2925 1078 2959 1112
rect 2993 1078 3027 1112
rect 3061 1078 3095 1112
rect 3129 1078 3163 1112
rect 3197 1078 3231 1112
rect 3265 1078 3299 1112
rect 3333 1078 3367 1112
rect 3401 1078 3435 1112
rect -10 986 24 1020
rect -10 918 24 952
rect -10 850 24 884
rect -10 782 24 816
rect -10 714 24 748
rect -10 646 24 680
rect -10 578 24 612
rect -10 510 24 544
rect -10 442 24 476
rect -10 374 24 408
rect -10 306 24 340
rect -10 238 24 272
rect -10 170 24 204
rect -10 102 24 136
rect -10 34 24 68
rect -10 -34 24 0
rect 123 -150 157 -116
rect 191 -150 225 -116
rect 259 -150 293 -116
rect 327 -150 361 -116
rect 395 -150 429 -116
rect 463 -150 497 -116
rect 531 -150 565 -116
rect 599 -150 633 -116
rect 667 -150 701 -116
rect 735 -150 769 -116
rect 803 -150 837 -116
rect 871 -150 905 -116
rect 939 -150 973 -116
rect 1007 -150 1041 -116
rect 1075 -150 1109 -116
<< mvnsubdiffcont >>
rect 348 892 382 926
rect 416 892 450 926
rect 484 892 518 926
rect 655 892 689 926
rect 723 892 757 926
rect 791 892 825 926
rect 859 892 893 926
rect 927 892 961 926
rect 995 892 1029 926
rect 1063 892 1097 926
rect 1131 892 1165 926
rect 1199 892 1233 926
rect 1267 892 1301 926
rect 1335 892 1369 926
rect 1403 892 1437 926
rect 1471 892 1505 926
rect 1539 892 1573 926
rect 1607 892 1641 926
rect 1675 892 1709 926
rect 1743 892 1777 926
rect 1811 892 1845 926
rect 1879 892 1913 926
rect 1947 892 1981 926
rect 2015 892 2049 926
rect 2083 892 2117 926
rect 2151 892 2185 926
rect 2219 892 2253 926
rect 2287 892 2321 926
rect 2355 892 2389 926
rect 2423 892 2457 926
rect 2491 892 2525 926
rect 2559 892 2593 926
rect 2627 892 2661 926
rect 2695 892 2729 926
rect 2763 892 2797 926
rect 2831 892 2865 926
rect 2899 892 2933 926
rect 2967 892 3001 926
rect 3035 892 3069 926
rect 3103 892 3137 926
rect 3171 892 3205 926
rect 3239 892 3273 926
rect 3307 892 3341 926
rect 3375 892 3409 926
rect 324 808 358 842
rect 393 790 427 824
rect 467 790 501 824
rect 541 790 575 824
rect 3450 868 3484 902
rect 324 740 358 774
rect 3450 800 3484 834
rect 393 717 427 751
rect 467 717 501 751
rect 541 717 575 751
rect 324 672 358 706
rect 393 644 427 678
rect 467 644 501 678
rect 541 644 575 678
rect 324 604 358 638
rect 393 571 427 605
rect 467 571 501 605
rect 541 571 575 605
rect 324 536 358 570
rect 324 468 358 502
rect 393 498 427 532
rect 467 498 501 532
rect 541 498 575 532
rect 324 400 358 434
rect 393 425 427 459
rect 467 425 501 459
rect 541 425 575 459
rect 324 332 358 366
rect 393 352 427 386
rect 467 352 501 386
rect 541 352 575 386
rect 324 264 358 298
rect 393 278 427 312
rect 467 278 501 312
rect 541 278 575 312
rect 324 196 358 230
rect 393 204 427 238
rect 467 204 501 238
rect 541 204 575 238
rect 3450 732 3484 766
rect 3450 664 3484 698
rect 3450 596 3484 630
rect 3450 528 3484 562
rect 3450 460 3484 494
rect 3450 392 3484 426
rect 3450 324 3484 358
rect 3450 256 3484 290
rect 324 128 358 162
rect 393 130 427 164
rect 467 130 501 164
rect 541 130 575 164
rect 3450 188 3484 222
rect 324 60 358 94
rect 3450 120 3484 154
rect 434 36 468 70
rect 502 36 536 70
rect 570 36 604 70
rect 638 36 672 70
rect 706 36 740 70
rect 774 36 808 70
rect 842 36 876 70
rect 910 36 944 70
rect 978 36 1012 70
rect 1046 36 1080 70
rect 1114 36 1148 70
rect 1182 36 1216 70
rect 1250 36 1284 70
rect 1318 36 1352 70
rect 1386 36 1420 70
rect 1454 36 1488 70
rect 1522 36 1556 70
rect 1590 36 1624 70
rect 1658 36 1692 70
rect 1726 36 1760 70
rect 1794 36 1828 70
rect 1862 36 1896 70
rect 1930 36 1964 70
rect 1998 36 2032 70
rect 2066 36 2100 70
rect 2134 36 2168 70
rect 2202 36 2236 70
rect 2270 36 2304 70
rect 2338 36 2372 70
rect 2406 36 2440 70
rect 2474 36 2508 70
rect 2542 36 2576 70
rect 2610 36 2644 70
rect 2678 36 2712 70
rect 2746 36 2780 70
rect 2814 36 2848 70
rect 2882 36 2916 70
rect 2950 36 2984 70
rect 3018 36 3052 70
rect 3086 36 3120 70
rect 3154 36 3188 70
rect 3222 36 3256 70
rect 3290 36 3324 70
rect 3358 36 3392 70
rect 3426 36 3460 70
<< poly >>
rect 652 749 756 765
rect 652 715 674 749
rect 708 715 756 749
rect 652 677 756 715
rect 652 643 674 677
rect 708 665 756 677
rect 1756 746 1886 765
rect 1756 712 1804 746
rect 1838 712 1886 746
rect 1756 674 1886 712
rect 1756 665 1804 674
rect 708 643 730 665
rect 652 609 730 643
rect 1782 640 1804 665
rect 1838 665 1886 674
rect 3286 746 3390 765
rect 3286 712 3334 746
rect 3368 712 3390 746
rect 3286 674 3390 712
rect 3286 665 3334 674
rect 1838 640 1860 665
rect 1782 609 1860 640
rect 3312 640 3334 665
rect 3368 640 3390 674
rect 3312 609 3390 640
rect 652 605 756 609
rect 652 571 674 605
rect 708 571 756 605
rect 652 533 756 571
rect 652 499 674 533
rect 708 509 756 533
rect 1756 602 1886 609
rect 1756 568 1804 602
rect 1838 568 1886 602
rect 1756 531 1886 568
rect 1756 509 1804 531
rect 708 499 730 509
rect 652 461 730 499
rect 652 427 674 461
rect 708 453 730 461
rect 1782 497 1804 509
rect 1838 509 1886 531
rect 3286 602 3390 609
rect 3286 568 3334 602
rect 3368 568 3390 602
rect 3286 531 3390 568
rect 3286 509 3334 531
rect 1838 497 1860 509
rect 1782 460 1860 497
rect 1782 453 1804 460
rect 708 427 756 453
rect 652 389 756 427
rect 652 355 674 389
rect 708 355 756 389
rect 652 353 756 355
rect 1756 426 1804 453
rect 1838 453 1860 460
rect 3312 497 3334 509
rect 3368 497 3390 531
rect 3312 460 3390 497
rect 3312 453 3334 460
rect 1838 426 1886 453
rect 1756 389 1886 426
rect 1756 355 1804 389
rect 1838 355 1886 389
rect 1756 353 1886 355
rect 3286 426 3334 453
rect 3368 426 3390 460
rect 3286 389 3390 426
rect 3286 355 3334 389
rect 3368 355 3390 389
rect 3286 353 3390 355
rect 652 318 730 353
rect 652 284 674 318
rect 708 297 730 318
rect 1782 318 1860 353
rect 1782 297 1804 318
rect 708 284 756 297
rect 652 247 756 284
rect 652 213 674 247
rect 708 213 756 247
rect 652 197 756 213
rect 1756 284 1804 297
rect 1838 297 1860 318
rect 3312 318 3390 353
rect 3312 297 3334 318
rect 1838 284 1886 297
rect 1756 247 1886 284
rect 1756 213 1804 247
rect 1838 213 1886 247
rect 1756 197 1886 213
rect 3286 284 3334 297
rect 3368 284 3390 318
rect 3286 247 3390 284
rect 3286 213 3334 247
rect 3368 213 3390 247
rect 3286 197 3390 213
<< polycont >>
rect 674 715 708 749
rect 674 643 708 677
rect 1804 712 1838 746
rect 1804 640 1838 674
rect 3334 712 3368 746
rect 3334 640 3368 674
rect 674 571 708 605
rect 674 499 708 533
rect 1804 568 1838 602
rect 674 427 708 461
rect 1804 497 1838 531
rect 3334 568 3368 602
rect 674 355 708 389
rect 1804 426 1838 460
rect 3334 497 3368 531
rect 1804 355 1838 389
rect 3334 426 3368 460
rect 3334 355 3368 389
rect 674 284 708 318
rect 674 213 708 247
rect 1804 284 1838 318
rect 1804 213 1838 247
rect 3334 284 3368 318
rect 3334 213 3368 247
<< locali >>
rect -10 1100 69 1112
rect 24 1078 69 1100
rect 135 1078 137 1112
rect 171 1078 173 1112
rect 239 1078 245 1112
rect 307 1078 317 1112
rect 375 1078 389 1112
rect 443 1078 461 1112
rect 511 1078 533 1112
rect 579 1078 605 1112
rect 647 1078 677 1112
rect 715 1078 749 1112
rect 783 1078 817 1112
rect 855 1078 885 1112
rect 927 1078 953 1112
rect 999 1078 1021 1112
rect 1071 1078 1089 1112
rect 1143 1078 1157 1112
rect 1215 1078 1225 1112
rect 1287 1078 1293 1112
rect 1359 1078 1361 1112
rect 1395 1078 1397 1112
rect 1463 1078 1469 1112
rect 1531 1078 1541 1112
rect 1599 1078 1613 1112
rect 1667 1078 1685 1112
rect 1735 1078 1757 1112
rect 1803 1078 1829 1112
rect 1871 1078 1901 1112
rect 1939 1078 1973 1112
rect 2007 1078 2041 1112
rect 2079 1078 2109 1112
rect 2151 1078 2177 1112
rect 2223 1078 2245 1112
rect 2295 1078 2313 1112
rect 2367 1078 2381 1112
rect 2439 1078 2449 1112
rect 2511 1078 2517 1112
rect 2583 1078 2585 1112
rect 2619 1078 2621 1112
rect 2687 1078 2693 1112
rect 2755 1078 2765 1112
rect 2823 1078 2837 1112
rect 2891 1078 2909 1112
rect 2959 1078 2981 1112
rect 3027 1078 3053 1112
rect 3095 1078 3125 1112
rect 3163 1078 3197 1112
rect 3231 1078 3265 1112
rect 3303 1078 3333 1112
rect 3375 1078 3401 1112
rect 3447 1078 3475 1112
rect -10 1028 24 1054
rect -10 956 24 986
rect -10 884 24 918
rect -10 816 24 850
rect -10 748 24 778
rect -10 680 24 706
rect -10 612 24 634
rect -10 544 24 562
rect -10 476 24 490
rect -10 408 24 418
rect -10 340 24 346
rect -10 272 24 274
rect -10 236 24 238
rect -10 164 24 170
rect -10 92 24 102
rect 324 892 336 926
rect 382 892 408 926
rect 450 892 480 926
rect 518 892 655 926
rect 689 892 723 926
rect 761 892 791 926
rect 833 892 859 926
rect 905 892 927 926
rect 977 892 995 926
rect 1049 892 1063 926
rect 1121 892 1131 926
rect 1193 892 1199 926
rect 1265 892 1267 926
rect 1301 892 1303 926
rect 1369 892 1375 926
rect 1437 892 1447 926
rect 1505 892 1519 926
rect 1573 892 1591 926
rect 1641 892 1663 926
rect 1709 892 1735 926
rect 1777 892 1807 926
rect 1845 892 1879 926
rect 1913 892 1947 926
rect 1985 892 2015 926
rect 2057 892 2083 926
rect 2129 892 2151 926
rect 2201 892 2219 926
rect 2273 892 2287 926
rect 2321 892 2355 926
rect 2389 892 2423 926
rect 2457 892 2491 926
rect 2525 892 2559 926
rect 2593 892 2627 926
rect 2661 892 2695 926
rect 2729 892 2763 926
rect 2797 892 2831 926
rect 2865 892 2899 926
rect 2933 892 2967 926
rect 3001 892 3035 926
rect 3069 892 3103 926
rect 3137 892 3171 926
rect 3205 892 3239 926
rect 3273 892 3307 926
rect 3341 892 3375 926
rect 3409 902 3484 926
rect 3409 892 3450 902
rect 324 842 575 892
rect 358 824 575 842
rect 358 808 393 824
rect 427 821 467 824
rect 324 802 393 808
rect 358 790 393 802
rect 459 790 467 821
rect 501 821 541 824
rect 501 790 529 821
rect 3450 834 3484 868
rect 358 787 425 790
rect 459 787 529 790
rect 563 787 575 790
rect 358 751 575 787
rect 824 776 826 810
rect 860 776 862 810
rect 928 776 934 810
rect 996 776 1006 810
rect 1064 776 1078 810
rect 1132 776 1150 810
rect 1200 776 1222 810
rect 1268 776 1294 810
rect 1336 776 1366 810
rect 1404 776 1438 810
rect 1472 776 1506 810
rect 1544 776 1574 810
rect 1616 776 1642 810
rect 1688 776 1710 810
rect 1922 776 1948 810
rect 1994 776 2016 810
rect 2066 776 2084 810
rect 2138 776 2152 810
rect 2210 776 2220 810
rect 2282 776 2288 810
rect 2354 776 2356 810
rect 2390 776 2392 810
rect 2458 776 2464 810
rect 2526 776 2536 810
rect 2594 776 2608 810
rect 2662 776 2680 810
rect 2730 776 2752 810
rect 2798 776 2824 810
rect 2866 776 2896 810
rect 2934 776 2968 810
rect 3002 776 3036 810
rect 3074 776 3104 810
rect 3146 776 3172 810
rect 3218 776 3240 810
rect 3450 766 3484 800
rect 358 740 393 751
rect 324 730 393 740
rect 358 717 393 730
rect 427 717 467 751
rect 501 717 541 751
rect 358 678 575 717
rect 358 672 393 678
rect 324 658 393 672
rect 358 644 393 658
rect 427 644 467 678
rect 501 644 541 678
rect 358 605 575 644
rect 358 604 393 605
rect 324 586 393 604
rect 358 571 393 586
rect 427 571 467 605
rect 501 571 541 605
rect 358 536 575 571
rect 324 532 575 536
rect 324 514 393 532
rect 358 498 393 514
rect 427 498 467 532
rect 501 498 541 532
rect 358 468 575 498
rect 324 459 575 468
rect 324 442 393 459
rect 358 425 393 442
rect 427 425 467 459
rect 501 425 541 459
rect 358 400 575 425
rect 324 386 575 400
rect 324 370 393 386
rect 358 352 393 370
rect 427 352 467 386
rect 501 352 541 386
rect 358 332 575 352
rect 324 312 575 332
rect 324 298 393 312
rect 358 278 393 298
rect 427 278 467 312
rect 501 278 541 312
rect 358 264 575 278
rect 324 238 575 264
rect 324 230 393 238
rect 358 204 393 230
rect 427 204 467 238
rect 501 204 541 238
rect 358 192 575 204
rect 674 749 708 765
rect 674 677 708 715
rect 1804 746 1838 762
rect 1804 674 1838 712
rect 674 605 708 643
rect 824 620 826 654
rect 860 620 862 654
rect 928 620 934 654
rect 996 620 1006 654
rect 1064 620 1078 654
rect 1132 620 1150 654
rect 1200 620 1222 654
rect 1268 620 1294 654
rect 1336 620 1366 654
rect 1404 620 1438 654
rect 1472 620 1506 654
rect 1544 620 1574 654
rect 1616 620 1642 654
rect 1688 620 1710 654
rect 3334 746 3368 762
rect 3334 674 3368 712
rect 1804 602 1838 640
rect 1922 620 1948 654
rect 1994 620 2016 654
rect 2066 620 2084 654
rect 2138 620 2152 654
rect 2210 620 2220 654
rect 2282 620 2288 654
rect 2354 620 2356 654
rect 2390 620 2392 654
rect 2458 620 2464 654
rect 2526 620 2536 654
rect 2594 620 2608 654
rect 2662 620 2680 654
rect 2730 620 2752 654
rect 2798 620 2824 654
rect 2866 620 2896 654
rect 2934 620 2968 654
rect 3002 620 3036 654
rect 3074 620 3104 654
rect 3146 620 3172 654
rect 3218 620 3240 654
rect 3334 602 3368 640
rect 674 541 688 571
rect 722 541 760 575
rect 1838 568 1863 575
rect 1825 541 1863 568
rect 3295 541 3333 575
rect 3367 541 3368 568
rect 674 533 708 541
rect 674 461 708 499
rect 1804 531 1838 541
rect 824 464 826 498
rect 860 464 862 498
rect 928 464 934 498
rect 996 464 1006 498
rect 1064 464 1078 498
rect 1132 464 1150 498
rect 1200 464 1222 498
rect 1268 464 1294 498
rect 1336 464 1366 498
rect 1404 464 1438 498
rect 1472 464 1506 498
rect 1544 464 1574 498
rect 1616 464 1642 498
rect 1688 464 1710 498
rect 3334 531 3368 541
rect 674 389 708 427
rect 674 318 708 355
rect 1804 460 1838 497
rect 1922 464 1948 498
rect 1994 464 2016 498
rect 2066 464 2084 498
rect 2138 464 2152 498
rect 2210 464 2220 498
rect 2282 464 2288 498
rect 2354 464 2356 498
rect 2390 464 2392 498
rect 2458 464 2464 498
rect 2526 464 2536 498
rect 2594 464 2608 498
rect 2662 464 2680 498
rect 2730 464 2752 498
rect 2798 464 2824 498
rect 2866 464 2896 498
rect 2934 464 2968 498
rect 3002 464 3036 498
rect 3074 464 3104 498
rect 3146 464 3172 498
rect 3218 464 3240 498
rect 1804 389 1838 426
rect 824 308 826 342
rect 860 308 862 342
rect 928 308 934 342
rect 996 308 1006 342
rect 1064 308 1078 342
rect 1132 308 1150 342
rect 1200 308 1222 342
rect 1268 308 1294 342
rect 1336 308 1366 342
rect 1404 308 1438 342
rect 1472 308 1506 342
rect 1544 308 1574 342
rect 1616 308 1642 342
rect 1688 308 1710 342
rect 1804 318 1838 355
rect 3334 460 3368 497
rect 3334 389 3368 426
rect 674 247 708 284
rect 674 197 708 213
rect 1922 308 1948 342
rect 1994 308 2016 342
rect 2066 308 2084 342
rect 2138 308 2152 342
rect 2210 308 2220 342
rect 2282 308 2288 342
rect 2354 308 2356 342
rect 2390 308 2392 342
rect 2458 308 2464 342
rect 2526 308 2536 342
rect 2594 308 2608 342
rect 2662 308 2680 342
rect 2730 308 2752 342
rect 2798 308 2824 342
rect 2866 308 2896 342
rect 2934 308 2968 342
rect 3002 308 3036 342
rect 3074 308 3104 342
rect 3146 308 3172 342
rect 3218 308 3240 342
rect 3334 318 3368 355
rect 1804 247 1838 284
rect 1804 197 1838 213
rect 3334 247 3368 284
rect 3334 197 3368 213
rect 3450 698 3484 732
rect 3450 630 3484 664
rect 3450 562 3484 596
rect 3450 494 3484 528
rect 3450 426 3484 460
rect 3450 358 3484 392
rect 3450 290 3484 324
rect 3450 222 3484 256
rect 324 179 575 192
rect 324 164 425 179
rect 459 164 529 179
rect 563 164 575 179
rect 324 162 393 164
rect 358 130 393 162
rect 459 145 467 164
rect 427 130 467 145
rect 501 145 529 164
rect 824 152 826 186
rect 860 152 862 186
rect 928 152 934 186
rect 996 152 1006 186
rect 1064 152 1078 186
rect 1132 152 1150 186
rect 1200 152 1222 186
rect 1268 152 1294 186
rect 1336 152 1366 186
rect 1404 152 1438 186
rect 1472 152 1506 186
rect 1544 152 1574 186
rect 1616 152 1642 186
rect 1688 152 1710 186
rect 1922 152 1948 186
rect 1994 152 2016 186
rect 2066 152 2084 186
rect 2138 152 2152 186
rect 2210 152 2220 186
rect 2282 152 2288 186
rect 2354 152 2356 186
rect 2390 152 2392 186
rect 2458 152 2464 186
rect 2526 152 2536 186
rect 2594 152 2608 186
rect 2662 152 2680 186
rect 2730 152 2752 186
rect 2798 152 2824 186
rect 2866 152 2896 186
rect 2934 152 2968 186
rect 3002 152 3036 186
rect 3074 152 3104 186
rect 3146 152 3172 186
rect 3218 152 3240 186
rect 3450 154 3484 188
rect 501 130 541 145
rect 358 120 575 130
rect 324 94 575 120
rect 358 70 575 94
rect 3450 70 3484 120
rect 358 48 434 70
rect 324 36 434 48
rect 500 36 502 70
rect 536 36 538 70
rect 604 36 610 70
rect 672 36 682 70
rect 740 36 754 70
rect 808 36 826 70
rect 876 36 898 70
rect 944 36 970 70
rect 1012 36 1042 70
rect 1080 36 1114 70
rect 1148 36 1182 70
rect 1220 36 1250 70
rect 1292 36 1318 70
rect 1364 36 1386 70
rect 1436 36 1454 70
rect 1508 36 1522 70
rect 1580 36 1590 70
rect 1652 36 1658 70
rect 1724 36 1726 70
rect 1760 36 1762 70
rect 1828 36 1834 70
rect 1896 36 1906 70
rect 1964 36 1978 70
rect 2032 36 2050 70
rect 2100 36 2122 70
rect 2168 36 2194 70
rect 2236 36 2266 70
rect 2304 36 2338 70
rect 2372 36 2406 70
rect 2444 36 2474 70
rect 2516 36 2542 70
rect 2588 36 2610 70
rect 2660 36 2678 70
rect 2732 36 2746 70
rect 2804 36 2814 70
rect 2876 36 2882 70
rect 2948 36 2950 70
rect 2984 36 2986 70
rect 3052 36 3058 70
rect 3120 36 3130 70
rect 3188 36 3202 70
rect 3256 36 3274 70
rect 3324 36 3346 70
rect 3392 36 3426 70
rect 3460 36 3484 70
rect -10 20 24 34
rect -10 -116 24 -34
rect -10 -150 111 -116
rect 157 -150 183 -116
rect 225 -150 255 -116
rect 293 -150 327 -116
rect 361 -150 395 -116
rect 433 -150 463 -116
rect 505 -150 531 -116
rect 577 -150 599 -116
rect 649 -150 667 -116
rect 721 -150 735 -116
rect 793 -150 803 -116
rect 865 -150 871 -116
rect 937 -150 939 -116
rect 973 -150 975 -116
rect 1041 -150 1047 -116
rect 1109 -150 1119 -116
rect 1153 -138 1193 -116
rect 1227 -138 1266 -104
rect 1300 -138 1339 -104
rect 1373 -138 1412 -104
rect 1446 -138 1485 -104
rect 1519 -138 1558 -104
rect 1592 -138 1631 -104
rect 1665 -138 1704 -104
rect 1738 -138 1777 -104
rect 1811 -138 1850 -104
rect 1884 -138 1923 -104
rect 1957 -138 1996 -104
rect 2030 -138 2069 -104
rect 2103 -138 2142 -104
rect 2176 -138 2216 -104
rect 2250 -138 2290 -104
rect 2324 -138 2364 -104
rect 2398 -138 2438 -104
rect 2472 -138 2512 -104
rect 2546 -138 2586 -104
rect 2620 -138 2660 -104
rect 2694 -138 2734 -104
rect 2768 -138 2808 -104
rect 2842 -138 2882 -104
rect 2916 -138 2956 -104
rect 2990 -138 3030 -104
rect 3064 -138 3104 -104
rect 3138 -138 3178 -104
rect 3212 -138 3252 -104
rect 3286 -138 3326 -104
rect 3360 -138 3400 -104
rect 3434 -138 3467 -116
rect 1153 -150 3467 -138
<< viali >>
rect -10 1088 24 1100
rect -10 1066 24 1088
rect 101 1078 103 1112
rect 103 1078 135 1112
rect 173 1078 205 1112
rect 205 1078 207 1112
rect 245 1078 273 1112
rect 273 1078 279 1112
rect 317 1078 341 1112
rect 341 1078 351 1112
rect 389 1078 409 1112
rect 409 1078 423 1112
rect 461 1078 477 1112
rect 477 1078 495 1112
rect 533 1078 545 1112
rect 545 1078 567 1112
rect 605 1078 613 1112
rect 613 1078 639 1112
rect 677 1078 681 1112
rect 681 1078 711 1112
rect 749 1078 783 1112
rect 821 1078 851 1112
rect 851 1078 855 1112
rect 893 1078 919 1112
rect 919 1078 927 1112
rect 965 1078 987 1112
rect 987 1078 999 1112
rect 1037 1078 1055 1112
rect 1055 1078 1071 1112
rect 1109 1078 1123 1112
rect 1123 1078 1143 1112
rect 1181 1078 1191 1112
rect 1191 1078 1215 1112
rect 1253 1078 1259 1112
rect 1259 1078 1287 1112
rect 1325 1078 1327 1112
rect 1327 1078 1359 1112
rect 1397 1078 1429 1112
rect 1429 1078 1431 1112
rect 1469 1078 1497 1112
rect 1497 1078 1503 1112
rect 1541 1078 1565 1112
rect 1565 1078 1575 1112
rect 1613 1078 1633 1112
rect 1633 1078 1647 1112
rect 1685 1078 1701 1112
rect 1701 1078 1719 1112
rect 1757 1078 1769 1112
rect 1769 1078 1791 1112
rect 1829 1078 1837 1112
rect 1837 1078 1863 1112
rect 1901 1078 1905 1112
rect 1905 1078 1935 1112
rect 1973 1078 2007 1112
rect 2045 1078 2075 1112
rect 2075 1078 2079 1112
rect 2117 1078 2143 1112
rect 2143 1078 2151 1112
rect 2189 1078 2211 1112
rect 2211 1078 2223 1112
rect 2261 1078 2279 1112
rect 2279 1078 2295 1112
rect 2333 1078 2347 1112
rect 2347 1078 2367 1112
rect 2405 1078 2415 1112
rect 2415 1078 2439 1112
rect 2477 1078 2483 1112
rect 2483 1078 2511 1112
rect 2549 1078 2551 1112
rect 2551 1078 2583 1112
rect 2621 1078 2653 1112
rect 2653 1078 2655 1112
rect 2693 1078 2721 1112
rect 2721 1078 2727 1112
rect 2765 1078 2789 1112
rect 2789 1078 2799 1112
rect 2837 1078 2857 1112
rect 2857 1078 2871 1112
rect 2909 1078 2925 1112
rect 2925 1078 2943 1112
rect 2981 1078 2993 1112
rect 2993 1078 3015 1112
rect 3053 1078 3061 1112
rect 3061 1078 3087 1112
rect 3125 1078 3129 1112
rect 3129 1078 3159 1112
rect 3197 1078 3231 1112
rect 3269 1078 3299 1112
rect 3299 1078 3303 1112
rect 3341 1078 3367 1112
rect 3367 1078 3375 1112
rect 3413 1078 3435 1112
rect 3435 1078 3447 1112
rect -10 1020 24 1028
rect -10 994 24 1020
rect -10 952 24 956
rect -10 922 24 952
rect -10 850 24 884
rect -10 782 24 812
rect -10 778 24 782
rect -10 714 24 740
rect -10 706 24 714
rect -10 646 24 668
rect -10 634 24 646
rect -10 578 24 596
rect -10 562 24 578
rect -10 510 24 524
rect -10 490 24 510
rect -10 442 24 452
rect -10 418 24 442
rect -10 374 24 380
rect -10 346 24 374
rect -10 306 24 308
rect -10 274 24 306
rect -10 204 24 236
rect -10 202 24 204
rect -10 136 24 164
rect -10 130 24 136
rect -10 68 24 92
rect -10 58 24 68
rect 336 892 348 926
rect 348 892 370 926
rect 408 892 416 926
rect 416 892 442 926
rect 480 892 484 926
rect 484 892 514 926
rect 655 892 689 926
rect 727 892 757 926
rect 757 892 761 926
rect 799 892 825 926
rect 825 892 833 926
rect 871 892 893 926
rect 893 892 905 926
rect 943 892 961 926
rect 961 892 977 926
rect 1015 892 1029 926
rect 1029 892 1049 926
rect 1087 892 1097 926
rect 1097 892 1121 926
rect 1159 892 1165 926
rect 1165 892 1193 926
rect 1231 892 1233 926
rect 1233 892 1265 926
rect 1303 892 1335 926
rect 1335 892 1337 926
rect 1375 892 1403 926
rect 1403 892 1409 926
rect 1447 892 1471 926
rect 1471 892 1481 926
rect 1519 892 1539 926
rect 1539 892 1553 926
rect 1591 892 1607 926
rect 1607 892 1625 926
rect 1663 892 1675 926
rect 1675 892 1697 926
rect 1735 892 1743 926
rect 1743 892 1769 926
rect 1807 892 1811 926
rect 1811 892 1841 926
rect 1879 892 1913 926
rect 1951 892 1981 926
rect 1981 892 1985 926
rect 2023 892 2049 926
rect 2049 892 2057 926
rect 2095 892 2117 926
rect 2117 892 2129 926
rect 2167 892 2185 926
rect 2185 892 2201 926
rect 2239 892 2253 926
rect 2253 892 2273 926
rect 324 774 358 802
rect 425 790 427 821
rect 427 790 459 821
rect 529 790 541 821
rect 541 790 563 821
rect 425 787 459 790
rect 529 787 563 790
rect 324 768 358 774
rect 790 776 824 810
rect 862 776 894 810
rect 894 776 896 810
rect 934 776 962 810
rect 962 776 968 810
rect 1006 776 1030 810
rect 1030 776 1040 810
rect 1078 776 1098 810
rect 1098 776 1112 810
rect 1150 776 1166 810
rect 1166 776 1184 810
rect 1222 776 1234 810
rect 1234 776 1256 810
rect 1294 776 1302 810
rect 1302 776 1328 810
rect 1366 776 1370 810
rect 1370 776 1400 810
rect 1438 776 1472 810
rect 1510 776 1540 810
rect 1540 776 1544 810
rect 1582 776 1608 810
rect 1608 776 1616 810
rect 1654 776 1676 810
rect 1676 776 1688 810
rect 1726 776 1744 810
rect 1744 776 1760 810
rect 1888 776 1922 810
rect 1960 776 1982 810
rect 1982 776 1994 810
rect 2032 776 2050 810
rect 2050 776 2066 810
rect 2104 776 2118 810
rect 2118 776 2138 810
rect 2176 776 2186 810
rect 2186 776 2210 810
rect 2248 776 2254 810
rect 2254 776 2282 810
rect 2320 776 2322 810
rect 2322 776 2354 810
rect 2392 776 2424 810
rect 2424 776 2426 810
rect 2464 776 2492 810
rect 2492 776 2498 810
rect 2536 776 2560 810
rect 2560 776 2570 810
rect 2608 776 2628 810
rect 2628 776 2642 810
rect 2680 776 2696 810
rect 2696 776 2714 810
rect 2752 776 2764 810
rect 2764 776 2786 810
rect 2824 776 2832 810
rect 2832 776 2858 810
rect 2896 776 2900 810
rect 2900 776 2930 810
rect 2968 776 3002 810
rect 3040 776 3070 810
rect 3070 776 3074 810
rect 3112 776 3138 810
rect 3138 776 3146 810
rect 3184 776 3206 810
rect 3206 776 3218 810
rect 3256 776 3274 810
rect 3274 776 3290 810
rect 324 706 358 730
rect 324 696 358 706
rect 324 638 358 658
rect 324 624 358 638
rect 324 570 358 586
rect 324 552 358 570
rect 324 502 358 514
rect 324 480 358 502
rect 324 434 358 442
rect 324 408 358 434
rect 324 366 358 370
rect 324 336 358 366
rect 324 264 358 298
rect 324 196 358 226
rect 324 192 358 196
rect 790 620 824 654
rect 862 620 894 654
rect 894 620 896 654
rect 934 620 962 654
rect 962 620 968 654
rect 1006 620 1030 654
rect 1030 620 1040 654
rect 1078 620 1098 654
rect 1098 620 1112 654
rect 1150 620 1166 654
rect 1166 620 1184 654
rect 1222 620 1234 654
rect 1234 620 1256 654
rect 1294 620 1302 654
rect 1302 620 1328 654
rect 1366 620 1370 654
rect 1370 620 1400 654
rect 1438 620 1472 654
rect 1510 620 1540 654
rect 1540 620 1544 654
rect 1582 620 1608 654
rect 1608 620 1616 654
rect 1654 620 1676 654
rect 1676 620 1688 654
rect 1726 620 1744 654
rect 1744 620 1760 654
rect 1888 620 1922 654
rect 1960 620 1982 654
rect 1982 620 1994 654
rect 2032 620 2050 654
rect 2050 620 2066 654
rect 2104 620 2118 654
rect 2118 620 2138 654
rect 2176 620 2186 654
rect 2186 620 2210 654
rect 2248 620 2254 654
rect 2254 620 2282 654
rect 2320 620 2322 654
rect 2322 620 2354 654
rect 2392 620 2424 654
rect 2424 620 2426 654
rect 2464 620 2492 654
rect 2492 620 2498 654
rect 2536 620 2560 654
rect 2560 620 2570 654
rect 2608 620 2628 654
rect 2628 620 2642 654
rect 2680 620 2696 654
rect 2696 620 2714 654
rect 2752 620 2764 654
rect 2764 620 2786 654
rect 2824 620 2832 654
rect 2832 620 2858 654
rect 2896 620 2900 654
rect 2900 620 2930 654
rect 2968 620 3002 654
rect 3040 620 3070 654
rect 3070 620 3074 654
rect 3112 620 3138 654
rect 3138 620 3146 654
rect 3184 620 3206 654
rect 3206 620 3218 654
rect 3256 620 3274 654
rect 3274 620 3290 654
rect 688 571 708 575
rect 708 571 722 575
rect 688 541 722 571
rect 760 541 794 575
rect 1791 568 1804 575
rect 1804 568 1825 575
rect 1791 541 1825 568
rect 1863 541 1897 575
rect 3261 541 3295 575
rect 3333 568 3334 575
rect 3334 568 3367 575
rect 3333 541 3367 568
rect 790 464 824 498
rect 862 464 894 498
rect 894 464 896 498
rect 934 464 962 498
rect 962 464 968 498
rect 1006 464 1030 498
rect 1030 464 1040 498
rect 1078 464 1098 498
rect 1098 464 1112 498
rect 1150 464 1166 498
rect 1166 464 1184 498
rect 1222 464 1234 498
rect 1234 464 1256 498
rect 1294 464 1302 498
rect 1302 464 1328 498
rect 1366 464 1370 498
rect 1370 464 1400 498
rect 1438 464 1472 498
rect 1510 464 1540 498
rect 1540 464 1544 498
rect 1582 464 1608 498
rect 1608 464 1616 498
rect 1654 464 1676 498
rect 1676 464 1688 498
rect 1726 464 1744 498
rect 1744 464 1760 498
rect 1888 464 1922 498
rect 1960 464 1982 498
rect 1982 464 1994 498
rect 2032 464 2050 498
rect 2050 464 2066 498
rect 2104 464 2118 498
rect 2118 464 2138 498
rect 2176 464 2186 498
rect 2186 464 2210 498
rect 2248 464 2254 498
rect 2254 464 2282 498
rect 2320 464 2322 498
rect 2322 464 2354 498
rect 2392 464 2424 498
rect 2424 464 2426 498
rect 2464 464 2492 498
rect 2492 464 2498 498
rect 2536 464 2560 498
rect 2560 464 2570 498
rect 2608 464 2628 498
rect 2628 464 2642 498
rect 2680 464 2696 498
rect 2696 464 2714 498
rect 2752 464 2764 498
rect 2764 464 2786 498
rect 2824 464 2832 498
rect 2832 464 2858 498
rect 2896 464 2900 498
rect 2900 464 2930 498
rect 2968 464 3002 498
rect 3040 464 3070 498
rect 3070 464 3074 498
rect 3112 464 3138 498
rect 3138 464 3146 498
rect 3184 464 3206 498
rect 3206 464 3218 498
rect 3256 464 3274 498
rect 3274 464 3290 498
rect 790 308 824 342
rect 862 308 894 342
rect 894 308 896 342
rect 934 308 962 342
rect 962 308 968 342
rect 1006 308 1030 342
rect 1030 308 1040 342
rect 1078 308 1098 342
rect 1098 308 1112 342
rect 1150 308 1166 342
rect 1166 308 1184 342
rect 1222 308 1234 342
rect 1234 308 1256 342
rect 1294 308 1302 342
rect 1302 308 1328 342
rect 1366 308 1370 342
rect 1370 308 1400 342
rect 1438 308 1472 342
rect 1510 308 1540 342
rect 1540 308 1544 342
rect 1582 308 1608 342
rect 1608 308 1616 342
rect 1654 308 1676 342
rect 1676 308 1688 342
rect 1726 308 1744 342
rect 1744 308 1760 342
rect 1888 308 1922 342
rect 1960 308 1982 342
rect 1982 308 1994 342
rect 2032 308 2050 342
rect 2050 308 2066 342
rect 2104 308 2118 342
rect 2118 308 2138 342
rect 2176 308 2186 342
rect 2186 308 2210 342
rect 2248 308 2254 342
rect 2254 308 2282 342
rect 2320 308 2322 342
rect 2322 308 2354 342
rect 2392 308 2424 342
rect 2424 308 2426 342
rect 2464 308 2492 342
rect 2492 308 2498 342
rect 2536 308 2560 342
rect 2560 308 2570 342
rect 2608 308 2628 342
rect 2628 308 2642 342
rect 2680 308 2696 342
rect 2696 308 2714 342
rect 2752 308 2764 342
rect 2764 308 2786 342
rect 2824 308 2832 342
rect 2832 308 2858 342
rect 2896 308 2900 342
rect 2900 308 2930 342
rect 2968 308 3002 342
rect 3040 308 3070 342
rect 3070 308 3074 342
rect 3112 308 3138 342
rect 3138 308 3146 342
rect 3184 308 3206 342
rect 3206 308 3218 342
rect 3256 308 3274 342
rect 3274 308 3290 342
rect 425 164 459 179
rect 529 164 563 179
rect 324 128 358 154
rect 425 145 427 164
rect 427 145 459 164
rect 529 145 541 164
rect 541 145 563 164
rect 790 152 824 186
rect 862 152 894 186
rect 894 152 896 186
rect 934 152 962 186
rect 962 152 968 186
rect 1006 152 1030 186
rect 1030 152 1040 186
rect 1078 152 1098 186
rect 1098 152 1112 186
rect 1150 152 1166 186
rect 1166 152 1184 186
rect 1222 152 1234 186
rect 1234 152 1256 186
rect 1294 152 1302 186
rect 1302 152 1328 186
rect 1366 152 1370 186
rect 1370 152 1400 186
rect 1438 152 1472 186
rect 1510 152 1540 186
rect 1540 152 1544 186
rect 1582 152 1608 186
rect 1608 152 1616 186
rect 1654 152 1676 186
rect 1676 152 1688 186
rect 1726 152 1744 186
rect 1744 152 1760 186
rect 1888 152 1922 186
rect 1960 152 1982 186
rect 1982 152 1994 186
rect 2032 152 2050 186
rect 2050 152 2066 186
rect 2104 152 2118 186
rect 2118 152 2138 186
rect 2176 152 2186 186
rect 2186 152 2210 186
rect 2248 152 2254 186
rect 2254 152 2282 186
rect 2320 152 2322 186
rect 2322 152 2354 186
rect 2392 152 2424 186
rect 2424 152 2426 186
rect 2464 152 2492 186
rect 2492 152 2498 186
rect 2536 152 2560 186
rect 2560 152 2570 186
rect 2608 152 2628 186
rect 2628 152 2642 186
rect 2680 152 2696 186
rect 2696 152 2714 186
rect 2752 152 2764 186
rect 2764 152 2786 186
rect 2824 152 2832 186
rect 2832 152 2858 186
rect 2896 152 2900 186
rect 2900 152 2930 186
rect 2968 152 3002 186
rect 3040 152 3070 186
rect 3070 152 3074 186
rect 3112 152 3138 186
rect 3138 152 3146 186
rect 3184 152 3206 186
rect 3206 152 3218 186
rect 3256 152 3274 186
rect 3274 152 3290 186
rect 324 120 358 128
rect 324 60 358 82
rect 324 48 358 60
rect 466 36 468 70
rect 468 36 500 70
rect 538 36 570 70
rect 570 36 572 70
rect 610 36 638 70
rect 638 36 644 70
rect 682 36 706 70
rect 706 36 716 70
rect 754 36 774 70
rect 774 36 788 70
rect 826 36 842 70
rect 842 36 860 70
rect 898 36 910 70
rect 910 36 932 70
rect 970 36 978 70
rect 978 36 1004 70
rect 1042 36 1046 70
rect 1046 36 1076 70
rect 1114 36 1148 70
rect 1186 36 1216 70
rect 1216 36 1220 70
rect 1258 36 1284 70
rect 1284 36 1292 70
rect 1330 36 1352 70
rect 1352 36 1364 70
rect 1402 36 1420 70
rect 1420 36 1436 70
rect 1474 36 1488 70
rect 1488 36 1508 70
rect 1546 36 1556 70
rect 1556 36 1580 70
rect 1618 36 1624 70
rect 1624 36 1652 70
rect 1690 36 1692 70
rect 1692 36 1724 70
rect 1762 36 1794 70
rect 1794 36 1796 70
rect 1834 36 1862 70
rect 1862 36 1868 70
rect 1906 36 1930 70
rect 1930 36 1940 70
rect 1978 36 1998 70
rect 1998 36 2012 70
rect 2050 36 2066 70
rect 2066 36 2084 70
rect 2122 36 2134 70
rect 2134 36 2156 70
rect 2194 36 2202 70
rect 2202 36 2228 70
rect 2266 36 2270 70
rect 2270 36 2300 70
rect 2338 36 2372 70
rect 2410 36 2440 70
rect 2440 36 2444 70
rect 2482 36 2508 70
rect 2508 36 2516 70
rect 2554 36 2576 70
rect 2576 36 2588 70
rect 2626 36 2644 70
rect 2644 36 2660 70
rect 2698 36 2712 70
rect 2712 36 2732 70
rect 2770 36 2780 70
rect 2780 36 2804 70
rect 2842 36 2848 70
rect 2848 36 2876 70
rect 2914 36 2916 70
rect 2916 36 2948 70
rect 2986 36 3018 70
rect 3018 36 3020 70
rect 3058 36 3086 70
rect 3086 36 3092 70
rect 3130 36 3154 70
rect 3154 36 3164 70
rect 3202 36 3222 70
rect 3222 36 3236 70
rect 3274 36 3290 70
rect 3290 36 3308 70
rect 3346 36 3358 70
rect 3358 36 3380 70
rect -10 0 24 20
rect -10 -14 24 0
rect 111 -150 123 -116
rect 123 -150 145 -116
rect 183 -150 191 -116
rect 191 -150 217 -116
rect 255 -150 259 -116
rect 259 -150 289 -116
rect 327 -150 361 -116
rect 399 -150 429 -116
rect 429 -150 433 -116
rect 471 -150 497 -116
rect 497 -150 505 -116
rect 543 -150 565 -116
rect 565 -150 577 -116
rect 615 -150 633 -116
rect 633 -150 649 -116
rect 687 -150 701 -116
rect 701 -150 721 -116
rect 759 -150 769 -116
rect 769 -150 793 -116
rect 831 -150 837 -116
rect 837 -150 865 -116
rect 903 -150 905 -116
rect 905 -150 937 -116
rect 975 -150 1007 -116
rect 1007 -150 1009 -116
rect 1047 -150 1075 -116
rect 1075 -150 1081 -116
rect 1119 -150 1153 -116
rect 1193 -138 1227 -104
rect 1266 -138 1300 -104
rect 1339 -138 1373 -104
rect 1412 -138 1446 -104
rect 1485 -138 1519 -104
rect 1558 -138 1592 -104
rect 1631 -138 1665 -104
rect 1704 -138 1738 -104
rect 1777 -138 1811 -104
rect 1850 -138 1884 -104
rect 1923 -138 1957 -104
rect 1996 -138 2030 -104
rect 2069 -138 2103 -104
rect 2142 -138 2176 -104
rect 2216 -138 2250 -104
rect 2290 -138 2324 -104
rect 2364 -138 2398 -104
rect 2438 -138 2472 -104
rect 2512 -138 2546 -104
rect 2586 -138 2620 -104
rect 2660 -138 2694 -104
rect 2734 -138 2768 -104
rect 2808 -138 2842 -104
rect 2882 -138 2916 -104
rect 2956 -138 2990 -104
rect 3030 -138 3064 -104
rect 3104 -138 3138 -104
rect 3178 -138 3212 -104
rect 3252 -138 3286 -104
rect 3326 -138 3360 -104
rect 3400 -138 3434 -104
<< metal1 >>
rect -22 1112 3467 1143
rect -22 1100 101 1112
rect -22 1066 -10 1100
rect 24 1078 101 1100
rect 135 1078 173 1112
rect 207 1078 245 1112
rect 279 1078 317 1112
rect 351 1078 389 1112
rect 423 1078 461 1112
rect 495 1078 533 1112
rect 567 1078 605 1112
rect 639 1078 677 1112
rect 711 1078 749 1112
rect 783 1078 821 1112
rect 855 1078 893 1112
rect 927 1078 965 1112
rect 999 1078 1037 1112
rect 1071 1078 1109 1112
rect 1143 1078 1181 1112
rect 1215 1078 1253 1112
rect 1287 1078 1325 1112
rect 1359 1078 1397 1112
rect 1431 1078 1469 1112
rect 1503 1078 1541 1112
rect 1575 1078 1613 1112
rect 1647 1078 1685 1112
rect 1719 1078 1757 1112
rect 1791 1078 1829 1112
rect 1863 1078 1901 1112
rect 1935 1078 1973 1112
rect 2007 1078 2045 1112
rect 2079 1078 2117 1112
rect 2151 1078 2189 1112
rect 2223 1078 2261 1112
rect 2295 1078 2333 1112
rect 2367 1078 2405 1112
rect 2439 1078 2477 1112
rect 2511 1078 2549 1112
rect 2583 1078 2621 1112
rect 2655 1078 2693 1112
rect 2727 1078 2765 1112
rect 2799 1078 2837 1112
rect 2871 1078 2909 1112
rect 2943 1078 2981 1112
rect 3015 1078 3053 1112
rect 3087 1078 3125 1112
rect 3159 1078 3197 1112
rect 3231 1078 3269 1112
rect 3303 1078 3341 1112
rect 3375 1078 3413 1112
rect 3447 1078 3467 1112
rect 24 1066 3467 1078
rect -22 1028 44 1066
rect -22 994 -10 1028
rect 24 994 44 1028
rect -22 956 44 994
rect -22 922 -10 956
rect 24 926 44 956
tri 44 926 184 1066 nw
rect 312 926 2370 938
rect 24 922 36 926
rect -22 884 36 922
tri 36 918 44 926 nw
rect -22 850 -10 884
rect 24 850 36 884
rect -22 812 36 850
rect -22 778 -10 812
rect 24 778 36 812
rect -22 740 36 778
rect -22 706 -10 740
rect 24 706 36 740
rect -22 668 36 706
rect -22 634 -10 668
rect 24 634 36 668
rect -22 596 36 634
rect -22 562 -10 596
rect 24 562 36 596
rect -22 524 36 562
rect -22 490 -10 524
rect 24 490 36 524
rect -22 452 36 490
rect -22 418 -10 452
rect 24 418 36 452
rect -22 380 36 418
rect -22 346 -10 380
rect 24 346 36 380
rect -22 308 36 346
rect -22 274 -10 308
rect 24 274 36 308
rect -22 236 36 274
rect -22 202 -10 236
rect 24 202 36 236
rect -22 164 36 202
rect -22 130 -10 164
rect 24 130 36 164
rect -22 92 36 130
rect -22 58 -10 92
rect 24 58 36 92
rect -22 36 36 58
rect 312 892 336 926
rect 370 892 408 926
rect 442 892 480 926
rect 514 892 655 926
rect 689 892 727 926
rect 761 892 799 926
rect 833 892 871 926
rect 905 892 943 926
rect 977 892 1015 926
rect 1049 892 1087 926
rect 1121 892 1159 926
rect 1193 892 1231 926
rect 1265 892 1303 926
rect 1337 892 1375 926
rect 1409 892 1447 926
rect 1481 892 1519 926
rect 1553 892 1591 926
rect 1625 892 1663 926
rect 1697 892 1735 926
rect 1769 892 1807 926
rect 1841 892 1879 926
rect 1913 892 1951 926
rect 1985 892 2023 926
rect 2057 892 2095 926
rect 2129 892 2167 926
rect 2201 892 2239 926
rect 2273 892 2370 926
rect 312 821 2370 892
rect 312 802 425 821
rect 312 768 324 802
rect 358 787 425 802
rect 459 787 529 821
rect 563 816 2370 821
rect 563 810 3496 816
rect 563 787 790 810
rect 358 776 790 787
rect 824 776 862 810
rect 896 776 934 810
rect 968 776 1006 810
rect 1040 776 1078 810
rect 1112 776 1150 810
rect 1184 776 1222 810
rect 1256 776 1294 810
rect 1328 776 1366 810
rect 1400 776 1438 810
rect 1472 776 1510 810
rect 1544 776 1582 810
rect 1616 776 1654 810
rect 1688 776 1726 810
rect 1760 776 1888 810
rect 1922 776 1960 810
rect 1994 776 2032 810
rect 2066 776 2104 810
rect 2138 776 2176 810
rect 2210 776 2248 810
rect 2282 776 2320 810
rect 2354 776 2392 810
rect 2426 776 2464 810
rect 2498 776 2536 810
rect 2570 776 2608 810
rect 2642 776 2680 810
rect 2714 776 2752 810
rect 2786 776 2824 810
rect 2858 776 2896 810
rect 2930 776 2968 810
rect 3002 776 3040 810
rect 3074 776 3112 810
rect 3146 776 3184 810
rect 3218 776 3256 810
rect 3290 805 3496 810
rect 3290 776 3438 805
rect 358 770 3438 776
rect 358 768 370 770
rect 312 730 370 768
tri 370 744 396 770 nw
tri 3379 744 3405 770 ne
rect 3405 744 3438 770
tri 3405 733 3416 744 ne
rect 3416 733 3438 744
rect 312 696 324 730
rect 358 696 370 730
rect 312 658 370 696
rect 312 624 324 658
rect 358 624 370 658
rect 312 586 370 624
rect 483 654 3302 733
tri 3416 711 3438 733 ne
rect 483 620 790 654
rect 824 620 862 654
rect 896 620 934 654
rect 968 620 1006 654
rect 1040 620 1078 654
rect 1112 620 1150 654
rect 1184 620 1222 654
rect 1256 620 1294 654
rect 1328 620 1366 654
rect 1400 620 1438 654
rect 1472 620 1510 654
rect 1544 620 1582 654
rect 1616 620 1654 654
rect 1688 620 1726 654
rect 1760 620 1888 654
rect 1922 620 1960 654
rect 1994 620 2032 654
rect 2066 620 2104 654
rect 2138 620 2176 654
rect 2210 620 2248 654
rect 2282 620 2320 654
rect 2354 620 2392 654
rect 2426 620 2464 654
rect 2498 620 2536 654
rect 2570 620 2608 654
rect 2642 620 2680 654
rect 2714 620 2752 654
rect 2786 620 2824 654
rect 2858 620 2896 654
rect 2930 620 2968 654
rect 3002 620 3040 654
rect 3074 620 3112 654
rect 3146 620 3184 654
rect 3218 620 3256 654
rect 3290 620 3302 654
rect 483 614 3302 620
rect 312 552 324 586
rect 358 552 370 586
rect 312 514 370 552
rect 676 575 3379 581
rect 676 541 688 575
rect 722 541 760 575
rect 794 541 1791 575
rect 1825 541 1863 575
rect 1897 541 3261 575
rect 3295 541 3333 575
rect 3367 541 3379 575
rect 676 535 3379 541
tri 3422 535 3438 551 se
tri 3420 533 3422 535 se
rect 3422 533 3438 535
rect 312 480 324 514
rect 358 504 370 514
tri 370 504 399 533 sw
tri 3391 504 3420 533 se
rect 3420 504 3438 533
rect 358 498 3438 504
rect 358 480 790 498
rect 312 464 790 480
rect 824 464 862 498
rect 896 464 934 498
rect 968 464 1006 498
rect 1040 464 1078 498
rect 1112 464 1150 498
rect 1184 464 1222 498
rect 1256 464 1294 498
rect 1328 464 1366 498
rect 1400 464 1438 498
rect 1472 464 1510 498
rect 1544 464 1582 498
rect 1616 464 1654 498
rect 1688 464 1726 498
rect 1760 464 1888 498
rect 1922 464 1960 498
rect 1994 464 2032 498
rect 2066 464 2104 498
rect 2138 464 2176 498
rect 2210 464 2248 498
rect 2282 464 2320 498
rect 2354 464 2392 498
rect 2426 464 2464 498
rect 2498 464 2536 498
rect 2570 464 2608 498
rect 2642 464 2680 498
rect 2714 464 2752 498
rect 2786 464 2824 498
rect 2858 464 2896 498
rect 2930 464 2968 498
rect 3002 464 3040 498
rect 3074 464 3112 498
rect 3146 464 3184 498
rect 3218 464 3256 498
rect 3290 464 3438 498
rect 312 442 3438 464
rect 312 408 324 442
rect 358 408 3438 442
rect 312 385 3438 408
rect 312 370 370 385
rect 312 336 324 370
rect 358 336 370 370
tri 370 354 401 385 nw
tri 3388 354 3419 385 ne
rect 3419 354 3438 385
tri 3419 348 3425 354 ne
rect 3425 348 3438 354
rect 312 298 370 336
rect 312 264 324 298
rect 358 264 370 298
rect 312 226 370 264
rect 407 342 3302 348
rect 407 308 790 342
rect 824 308 862 342
rect 896 308 934 342
rect 968 308 1006 342
rect 1040 308 1078 342
rect 1112 308 1150 342
rect 1184 308 1222 342
rect 1256 308 1294 342
rect 1328 308 1366 342
rect 1400 308 1438 342
rect 1472 308 1510 342
rect 1544 308 1582 342
rect 1616 308 1654 342
rect 1688 308 1726 342
rect 1760 308 1888 342
rect 1922 308 1960 342
rect 1994 308 2032 342
rect 2066 308 2104 342
rect 2138 308 2176 342
rect 2210 308 2248 342
rect 2282 308 2320 342
rect 2354 308 2392 342
rect 2426 308 2464 342
rect 2498 308 2536 342
rect 2570 308 2608 342
rect 2642 308 2680 342
rect 2714 308 2752 342
rect 2786 308 2824 342
rect 2858 308 2896 342
rect 2930 308 2968 342
rect 3002 308 3040 342
rect 3074 308 3112 342
rect 3146 308 3184 342
rect 3218 308 3256 342
rect 3290 308 3302 342
tri 3425 335 3438 348 ne
rect 407 279 3302 308
tri 407 229 457 279 ne
rect 457 229 3302 279
tri 3414 229 3444 259 se
rect 312 192 324 226
rect 358 192 370 226
tri 370 192 407 229 sw
tri 3377 192 3414 229 se
rect 3414 192 3444 229
rect 312 186 3444 192
rect 312 179 790 186
rect 312 154 425 179
rect 312 120 324 154
rect 358 145 425 154
rect 459 145 529 179
rect 563 152 790 179
rect 824 152 862 186
rect 896 152 934 186
rect 968 152 1006 186
rect 1040 152 1078 186
rect 1112 152 1150 186
rect 1184 152 1222 186
rect 1256 152 1294 186
rect 1328 152 1366 186
rect 1400 152 1438 186
rect 1472 152 1510 186
rect 1544 152 1582 186
rect 1616 152 1654 186
rect 1688 152 1726 186
rect 1760 152 1888 186
rect 1922 152 1960 186
rect 1994 152 2032 186
rect 2066 152 2104 186
rect 2138 152 2176 186
rect 2210 152 2248 186
rect 2282 152 2320 186
rect 2354 152 2392 186
rect 2426 152 2464 186
rect 2498 152 2536 186
rect 2570 152 2608 186
rect 2642 152 2680 186
rect 2714 152 2752 186
rect 2786 152 2824 186
rect 2858 152 2896 186
rect 2930 152 2968 186
rect 3002 152 3040 186
rect 3074 152 3112 186
rect 3146 152 3184 186
rect 3218 152 3256 186
rect 3290 152 3444 186
rect 563 145 3444 152
rect 358 120 3444 145
rect 312 104 3444 120
rect 312 89 3496 104
rect 312 82 3444 89
rect 312 48 324 82
rect 358 70 3444 82
rect 358 48 466 70
tri 36 36 38 38 sw
rect 312 36 466 48
rect 500 36 538 70
rect 572 36 610 70
rect 644 36 682 70
rect 716 36 754 70
rect 788 36 826 70
rect 860 36 898 70
rect 932 36 970 70
rect 1004 36 1042 70
rect 1076 36 1114 70
rect 1148 36 1186 70
rect 1220 36 1258 70
rect 1292 36 1330 70
rect 1364 36 1402 70
rect 1436 36 1474 70
rect 1508 36 1546 70
rect 1580 36 1618 70
rect 1652 36 1690 70
rect 1724 36 1762 70
rect 1796 36 1834 70
rect 1868 36 1906 70
rect 1940 36 1978 70
rect 2012 36 2050 70
rect 2084 36 2122 70
rect 2156 36 2194 70
rect 2228 36 2266 70
rect 2300 36 2338 70
rect 2372 36 2410 70
rect 2444 36 2482 70
rect 2516 36 2554 70
rect 2588 36 2626 70
rect 2660 36 2698 70
rect 2732 36 2770 70
rect 2804 36 2842 70
rect 2876 36 2914 70
rect 2948 36 2986 70
rect 3020 36 3058 70
rect 3092 36 3130 70
rect 3164 36 3202 70
rect 3236 36 3274 70
rect 3308 36 3346 70
rect 3380 67 3444 70
rect 3380 36 3420 67
rect -22 20 38 36
rect -22 -14 -10 20
rect 24 -14 38 20
rect -22 -70 38 -14
tri 38 -70 144 36 sw
rect 312 24 3420 36
rect -22 -104 144 -70
tri 144 -104 178 -70 sw
tri 1162 -104 1168 -98 se
rect 1168 -104 3488 -98
rect -22 -116 1193 -104
rect -22 -150 111 -116
rect 145 -150 183 -116
rect 217 -150 255 -116
rect 289 -150 327 -116
rect 361 -150 399 -116
rect 433 -150 471 -116
rect 505 -150 543 -116
rect 577 -150 615 -116
rect 649 -150 687 -116
rect 721 -150 759 -116
rect 793 -150 831 -116
rect 865 -150 903 -116
rect 937 -150 975 -116
rect 1009 -150 1047 -116
rect 1081 -150 1119 -116
rect 1153 -138 1193 -116
rect 1227 -138 1266 -104
rect 1300 -138 1339 -104
rect 1373 -138 1412 -104
rect 1446 -138 1485 -104
rect 1519 -138 1558 -104
rect 1592 -138 1631 -104
rect 1665 -138 1704 -104
rect 1738 -138 1777 -104
rect 1811 -138 1850 -104
rect 1884 -138 1923 -104
rect 1957 -138 1996 -104
rect 2030 -138 2069 -104
rect 2103 -138 2142 -104
rect 2176 -138 2216 -104
rect 2250 -138 2290 -104
rect 2324 -138 2364 -104
rect 2398 -138 2438 -104
rect 2472 -138 2512 -104
rect 2546 -138 2586 -104
rect 2620 -138 2660 -104
rect 2694 -138 2734 -104
rect 2768 -138 2808 -104
rect 2842 -138 2882 -104
rect 2916 -138 2956 -104
rect 2990 -138 3030 -104
rect 3064 -138 3104 -104
rect 3138 -138 3178 -104
rect 3212 -138 3252 -104
rect 3286 -138 3326 -104
rect 3360 -138 3400 -104
rect 3434 -138 3488 -104
rect 1153 -144 3488 -138
rect 1153 -150 1168 -144
rect -22 -162 1168 -150
tri 1168 -162 1186 -144 nw
use sky130_fd_pr__pfet_01v8__example_55959141808654  sky130_fd_pr__pfet_01v8__example_55959141808654_0
timestamp 1663361622
transform 0 -1 3286 1 0 197
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808656  sky130_fd_pr__pfet_01v8__example_55959141808656_0
timestamp 1663361622
transform 0 -1 1756 1 0 197
box -1 0 569 1
<< labels >>
flabel metal1 s 676 535 722 581 7 FreeSans 200 180 0 0 PU_H_N
port 1 nsew
flabel metal1 s 483 648 529 700 7 FreeSans 200 180 0 0 PAD
port 2 nsew
<< properties >>
string GDS_END 47424308
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 47390450
<< end >>
