magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 1 4 2 5 6 DRAIN
port 1 nsew
rlabel  s 1 5 2 5 6 DRAIN
port 1 nsew
rlabel  s 1 4 1 5 6 DRAIN
port 1 nsew
rlabel  s 0 5 2 6 6 GATE
port 2 nsew
rlabel  s 2 0 2 5 6 SOURCE
port 3 nsew
rlabel  s 1 0 1 5 6 SOURCE
port 3 nsew
rlabel  s 0 0 0 5 4 SOURCE
port 3 nsew
rlabel  s 0 0 2 0 8 SOURCE
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 2 6
string LEFview TRUE
<< end >>
