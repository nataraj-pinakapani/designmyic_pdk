magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 30 -17 64 21
<< locali >>
rect 103 333 169 493
rect 277 333 343 493
rect 103 299 359 333
rect 22 199 79 265
rect 119 199 195 265
rect 229 199 291 265
rect 119 60 162 199
rect 229 165 270 199
rect 325 165 359 299
rect 395 199 443 333
rect 200 60 270 165
rect 304 51 443 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 299 69 527
rect 203 367 237 527
rect 383 367 439 527
rect 18 17 85 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 395 199 443 333 6 A
port 1 nsew signal input
rlabel locali s 200 60 270 165 6 B
port 2 nsew signal input
rlabel locali s 229 165 270 199 6 B
port 2 nsew signal input
rlabel locali s 229 199 291 265 6 B
port 2 nsew signal input
rlabel locali s 119 60 162 199 6 C
port 3 nsew signal input
rlabel locali s 119 199 195 265 6 C
port 3 nsew signal input
rlabel locali s 22 199 79 265 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 459 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 304 51 443 165 6 Y
port 9 nsew signal output
rlabel locali s 325 165 359 299 6 Y
port 9 nsew signal output
rlabel locali s 103 299 359 333 6 Y
port 9 nsew signal output
rlabel locali s 277 333 343 493 6 Y
port 9 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1872856
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1867652
<< end >>
