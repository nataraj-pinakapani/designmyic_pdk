/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/openlane/custom_cells/lef/sky130_ef_io_core.lef