magic
tech sky130B
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__dfl1sd2__example_55959141808518  sky130_fd_pr__dfl1sd2__example_55959141808518_0
timestamp 1663361622
transform 1 0 160 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808517  sky130_fd_pr__dfl1sd__example_55959141808517_0
timestamp 1663361622
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808517  sky130_fd_pr__dfl1sd__example_55959141808517_1
timestamp 1663361622
transform 1 0 376 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 42393788
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 42392350
<< end >>
