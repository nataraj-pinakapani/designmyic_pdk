/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/ngspice/parasitics/sky130_fd_pr__model__parasitic__diodes_pw2dn.model.spice