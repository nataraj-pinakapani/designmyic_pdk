magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 46 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 54 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel 
 s 1 171 13 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel 
 s 1 24 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel 
 s 51 24 74 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel 
 s 62 171 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 198 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 13 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 174 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 51 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 198 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 62 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 198 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 197 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 197 75 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 75 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 75 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 75 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 195 75 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 195 75 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 75 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 75 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 75 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 193 75 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 193 75 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 75 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 75 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 75 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 191 75 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 191 75 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 75 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 75 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 75 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 189 75 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 189 75 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 75 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 75 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 75 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 187 75 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 187 75 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 75 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 75 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 75 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 185 75 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 185 75 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 75 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 75 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 75 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 183 75 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 183 75 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 75 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 75 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 75 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 181 75 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 181 75 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 75 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 75 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 75 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 179 75 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 179 75 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 75 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 75 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 75 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 177 75 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 177 75 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 75 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 75 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 75 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 175 75 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 175 75 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 174 75 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 174 75 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 198 74 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 197 74 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 197 74 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 74 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 74 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 74 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 195 74 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 195 74 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 74 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 74 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 74 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 193 74 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 193 74 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 74 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 74 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 74 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 191 74 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 191 74 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 74 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 74 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 74 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 189 74 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 189 74 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 74 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 74 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 74 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 187 74 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 187 74 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 74 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 74 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 74 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 185 74 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 185 74 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 74 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 74 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 74 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 183 74 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 183 74 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 74 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 74 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 74 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 181 74 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 181 74 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 74 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 74 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 74 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 179 74 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 179 74 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 74 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 74 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 74 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 177 74 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 177 74 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 74 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 74 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 74 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 175 74 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 175 74 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 174 74 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 174 74 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 28 74 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 28 74 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 27 74 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 27 74 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 26 74 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 26 74 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 26 74 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 25 74 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 25 74 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 24 74 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 24 74 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 198 74 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 197 74 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 197 74 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 74 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 74 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 196 74 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 195 74 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 195 74 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 74 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 74 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 194 74 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 193 74 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 193 74 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 74 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 74 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 192 74 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 191 74 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 191 74 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 74 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 74 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 190 74 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 189 74 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 189 74 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 74 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 74 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 188 74 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 187 74 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 187 74 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 74 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 74 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 186 74 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 185 74 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 185 74 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 74 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 74 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 184 74 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 183 74 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 183 74 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 74 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 74 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 182 74 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 181 74 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 181 74 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 74 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 74 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 180 74 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 179 74 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 179 74 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 74 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 74 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 178 74 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 177 74 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 177 74 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 74 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 74 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 176 74 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 175 74 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 175 74 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 174 74 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 174 74 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 28 74 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 28 74 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 27 74 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 27 74 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 26 74 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 26 74 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 26 74 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 25 74 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 25 74 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 24 74 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 74 24 74 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 198 73 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 197 73 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 197 73 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 196 73 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 196 73 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 196 73 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 195 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 195 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 194 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 194 73 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 194 73 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 193 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 193 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 192 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 192 73 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 192 73 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 191 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 191 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 190 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 190 73 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 190 73 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 189 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 189 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 188 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 188 73 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 188 73 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 187 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 187 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 186 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 186 73 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 186 73 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 185 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 185 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 184 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 184 73 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 184 73 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 183 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 183 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 182 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 182 73 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 182 73 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 181 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 181 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 180 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 180 73 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 180 73 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 179 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 179 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 178 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 178 73 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 178 73 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 177 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 177 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 176 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 176 73 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 176 73 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 175 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 175 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 174 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 174 73 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 28 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 28 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 27 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 27 73 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 26 73 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 26 73 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 26 73 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 25 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 25 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 24 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 24 73 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 198 73 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 197 73 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 197 73 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 196 73 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 196 73 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 196 73 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 195 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 195 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 194 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 194 73 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 194 73 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 193 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 193 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 192 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 192 73 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 192 73 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 191 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 191 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 190 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 190 73 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 190 73 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 189 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 189 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 188 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 188 73 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 188 73 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 187 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 187 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 186 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 186 73 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 186 73 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 185 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 185 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 184 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 184 73 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 184 73 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 183 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 183 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 182 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 182 73 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 182 73 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 181 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 181 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 180 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 180 73 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 180 73 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 179 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 179 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 178 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 178 73 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 178 73 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 177 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 177 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 176 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 176 73 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 176 73 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 175 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 175 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 174 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 174 73 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 28 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 28 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 27 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 27 73 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 26 73 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 26 73 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 26 73 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 25 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 25 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 24 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 73 24 73 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 198 73 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 197 73 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 197 73 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 73 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 73 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 73 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 195 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 195 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 73 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 73 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 73 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 193 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 193 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 73 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 73 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 73 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 191 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 191 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 73 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 73 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 73 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 189 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 189 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 73 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 73 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 73 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 187 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 187 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 73 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 73 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 73 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 185 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 185 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 73 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 73 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 73 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 183 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 183 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 73 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 73 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 73 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 181 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 181 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 73 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 73 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 73 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 179 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 179 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 73 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 73 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 73 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 177 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 177 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 73 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 73 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 73 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 175 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 175 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 174 73 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 174 73 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 28 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 28 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 27 73 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 27 73 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 73 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 73 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 73 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 25 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 25 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 24 73 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 24 73 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 198 72 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 197 72 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 197 72 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 72 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 72 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 72 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 195 72 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 195 72 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 72 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 72 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 72 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 193 72 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 193 72 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 72 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 72 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 72 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 191 72 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 191 72 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 72 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 72 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 72 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 189 72 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 189 72 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 72 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 72 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 72 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 187 72 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 187 72 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 72 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 72 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 72 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 185 72 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 185 72 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 72 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 72 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 72 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 183 72 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 183 72 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 72 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 72 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 72 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 181 72 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 181 72 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 72 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 72 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 72 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 179 72 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 179 72 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 72 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 72 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 72 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 177 72 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 177 72 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 72 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 72 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 72 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 175 72 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 175 72 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 174 72 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 174 72 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 28 72 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 28 72 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 27 72 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 27 72 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 72 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 72 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 72 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 25 72 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 25 72 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 24 72 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 24 72 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 198 72 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 197 72 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 197 72 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 72 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 72 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 196 72 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 195 72 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 195 72 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 72 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 72 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 194 72 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 193 72 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 193 72 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 72 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 72 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 192 72 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 191 72 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 191 72 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 72 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 72 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 190 72 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 189 72 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 189 72 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 72 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 72 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 188 72 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 187 72 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 187 72 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 72 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 72 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 186 72 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 185 72 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 185 72 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 72 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 72 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 184 72 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 183 72 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 183 72 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 72 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 72 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 182 72 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 181 72 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 181 72 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 72 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 72 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 180 72 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 179 72 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 179 72 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 72 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 72 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 178 72 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 177 72 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 177 72 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 72 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 72 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 176 72 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 175 72 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 175 72 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 174 72 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 174 72 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 28 72 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 28 72 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 27 72 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 27 72 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 72 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 72 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 26 72 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 25 72 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 25 72 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 24 72 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 72 24 72 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 28 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 28 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 27 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 27 71 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 26 71 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 26 71 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 26 71 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 25 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 25 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 24 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 24 71 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 198 71 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 197 71 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 197 71 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 196 71 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 196 71 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 196 71 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 195 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 195 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 194 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 194 71 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 194 71 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 193 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 193 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 192 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 192 71 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 192 71 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 191 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 191 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 190 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 190 71 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 190 71 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 189 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 189 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 188 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 188 71 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 188 71 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 187 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 187 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 186 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 186 71 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 186 71 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 185 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 185 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 184 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 184 71 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 184 71 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 183 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 183 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 182 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 182 71 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 182 71 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 181 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 181 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 180 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 180 71 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 180 71 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 179 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 179 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 178 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 178 71 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 178 71 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 177 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 177 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 176 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 176 71 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 176 71 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 175 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 175 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 174 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 174 71 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 28 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 28 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 27 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 27 71 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 26 71 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 26 71 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 26 71 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 25 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 25 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 24 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 24 71 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 198 71 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 197 71 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 197 71 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 196 71 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 196 71 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 196 71 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 195 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 195 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 194 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 194 71 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 194 71 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 193 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 193 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 192 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 192 71 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 192 71 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 191 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 191 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 190 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 190 71 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 190 71 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 189 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 189 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 188 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 188 71 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 188 71 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 187 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 187 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 186 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 186 71 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 186 71 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 185 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 185 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 184 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 184 71 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 184 71 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 183 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 183 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 182 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 182 71 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 182 71 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 181 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 181 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 180 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 180 71 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 180 71 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 179 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 179 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 178 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 178 71 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 178 71 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 177 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 177 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 176 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 176 71 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 176 71 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 175 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 175 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 174 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 71 174 71 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 28 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 28 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 27 71 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 27 71 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 71 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 71 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 71 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 25 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 25 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 24 71 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 24 71 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 198 71 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 197 71 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 197 71 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 71 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 71 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 71 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 195 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 195 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 71 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 71 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 71 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 193 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 193 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 71 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 71 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 71 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 191 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 191 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 71 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 71 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 71 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 189 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 189 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 71 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 71 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 71 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 187 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 187 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 71 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 71 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 71 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 185 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 185 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 71 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 71 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 71 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 183 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 183 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 71 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 71 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 71 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 181 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 181 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 71 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 71 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 71 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 179 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 179 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 71 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 71 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 71 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 177 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 177 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 71 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 71 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 71 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 175 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 175 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 174 71 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 174 71 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 28 70 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 28 70 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 27 70 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 27 70 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 70 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 70 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 70 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 25 70 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 25 70 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 24 70 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 24 70 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 198 70 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 197 70 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 197 70 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 70 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 70 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 70 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 195 70 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 195 70 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 70 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 70 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 70 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 193 70 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 193 70 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 70 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 70 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 70 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 191 70 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 191 70 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 70 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 70 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 70 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 189 70 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 189 70 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 70 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 70 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 70 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 187 70 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 187 70 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 70 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 70 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 70 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 185 70 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 185 70 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 70 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 70 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 70 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 183 70 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 183 70 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 70 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 70 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 70 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 181 70 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 181 70 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 70 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 70 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 70 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 179 70 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 179 70 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 70 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 70 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 70 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 177 70 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 177 70 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 70 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 70 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 70 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 175 70 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 175 70 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 174 70 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 174 70 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 28 70 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 28 70 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 27 70 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 27 70 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 70 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 70 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 26 70 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 25 70 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 25 70 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 24 70 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 24 70 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 198 70 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 197 70 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 197 70 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 70 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 70 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 196 70 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 195 70 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 195 70 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 70 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 70 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 194 70 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 193 70 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 193 70 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 70 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 70 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 192 70 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 191 70 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 191 70 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 70 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 70 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 190 70 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 189 70 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 189 70 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 70 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 70 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 188 70 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 187 70 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 187 70 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 70 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 70 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 186 70 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 185 70 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 185 70 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 70 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 70 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 184 70 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 183 70 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 183 70 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 70 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 70 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 182 70 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 181 70 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 181 70 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 70 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 70 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 180 70 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 179 70 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 179 70 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 70 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 70 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 178 70 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 177 70 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 177 70 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 70 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 70 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 176 70 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 175 70 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 175 70 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 174 70 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 70 174 70 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 28 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 28 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 27 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 27 69 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 26 69 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 26 69 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 26 69 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 25 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 25 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 24 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 24 69 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 198 69 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 197 69 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 197 69 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 196 69 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 196 69 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 196 69 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 195 69 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 195 69 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 194 69 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 194 69 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 194 69 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 193 69 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 193 69 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 192 69 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 192 69 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 192 69 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 191 69 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 191 69 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 190 69 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 190 69 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 190 69 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 189 69 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 189 69 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 188 69 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 188 69 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 188 69 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 187 69 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 187 69 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 186 69 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 186 69 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 186 69 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 185 69 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 185 69 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 184 69 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 184 69 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 184 69 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 183 69 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 183 69 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 182 69 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 182 69 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 182 69 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 181 69 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 181 69 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 180 69 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 180 69 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 180 69 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 179 69 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 179 69 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 178 69 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 178 69 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 178 69 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 177 69 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 177 69 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 176 69 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 176 69 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 176 69 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 175 69 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 175 69 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 174 69 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 174 69 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 28 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 28 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 27 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 27 69 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 26 69 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 26 69 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 26 69 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 25 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 25 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 24 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 24 69 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 198 69 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 197 69 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 197 69 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 196 69 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 196 69 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 196 69 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 195 69 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 195 69 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 194 69 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 194 69 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 194 69 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 193 69 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 193 69 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 192 69 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 192 69 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 192 69 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 191 69 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 191 69 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 190 69 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 190 69 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 190 69 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 189 69 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 189 69 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 188 69 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 188 69 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 188 69 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 187 69 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 187 69 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 186 69 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 186 69 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 186 69 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 185 69 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 185 69 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 184 69 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 184 69 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 184 69 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 183 69 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 183 69 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 182 69 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 182 69 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 182 69 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 181 69 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 181 69 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 180 69 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 180 69 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 180 69 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 179 69 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 179 69 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 178 69 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 178 69 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 178 69 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 177 69 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 177 69 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 176 69 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 176 69 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 176 69 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 175 69 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 175 69 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 174 69 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 69 174 69 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 28 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 28 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 27 69 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 27 69 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 69 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 69 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 69 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 25 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 25 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 24 69 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 24 69 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 198 68 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 197 68 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 197 68 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 196 68 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 196 68 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 196 68 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 195 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 195 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 194 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 194 68 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 194 68 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 193 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 193 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 192 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 192 68 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 192 68 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 191 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 191 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 190 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 190 68 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 190 68 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 189 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 189 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 188 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 188 68 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 188 68 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 187 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 187 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 186 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 186 68 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 186 68 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 185 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 185 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 184 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 184 68 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 184 68 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 183 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 183 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 182 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 182 68 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 182 68 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 181 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 181 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 180 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 180 68 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 180 68 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 179 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 179 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 178 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 178 68 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 178 68 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 177 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 177 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 176 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 176 68 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 176 68 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 175 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 175 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 174 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 174 68 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 28 68 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 28 68 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 27 68 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 27 68 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 68 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 68 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 68 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 25 68 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 25 68 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 24 68 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 24 68 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 198 68 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 197 68 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 197 68 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 196 68 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 196 68 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 196 68 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 195 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 195 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 194 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 194 68 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 194 68 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 193 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 193 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 192 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 192 68 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 192 68 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 191 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 191 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 190 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 190 68 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 190 68 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 189 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 189 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 188 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 188 68 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 188 68 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 187 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 187 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 186 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 186 68 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 186 68 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 185 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 185 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 184 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 184 68 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 184 68 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 183 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 183 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 182 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 182 68 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 182 68 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 181 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 181 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 180 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 180 68 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 180 68 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 179 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 179 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 178 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 178 68 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 178 68 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 177 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 177 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 176 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 176 68 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 176 68 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 175 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 175 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 174 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 174 68 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 28 68 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 28 68 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 27 68 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 27 68 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 68 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 68 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 26 68 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 25 68 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 25 68 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 24 68 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 68 24 68 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 198 68 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 197 68 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 197 68 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 68 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 68 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 68 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 195 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 195 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 68 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 68 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 68 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 193 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 193 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 68 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 68 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 68 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 191 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 191 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 68 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 68 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 68 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 189 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 189 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 68 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 68 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 68 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 187 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 187 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 68 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 68 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 68 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 185 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 185 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 68 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 68 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 68 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 183 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 183 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 68 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 68 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 68 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 181 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 181 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 68 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 68 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 68 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 179 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 179 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 68 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 68 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 68 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 177 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 177 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 68 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 68 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 68 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 175 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 175 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 174 68 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 174 68 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 28 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 28 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 27 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 27 67 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 26 67 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 26 67 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 26 67 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 25 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 25 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 24 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 24 67 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 198 67 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 197 67 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 197 67 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 67 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 67 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 67 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 195 67 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 195 67 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 67 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 67 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 67 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 193 67 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 193 67 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 67 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 67 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 67 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 191 67 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 191 67 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 67 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 67 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 67 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 189 67 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 189 67 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 67 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 67 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 67 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 187 67 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 187 67 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 67 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 67 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 67 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 185 67 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 185 67 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 67 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 67 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 67 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 183 67 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 183 67 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 67 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 67 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 67 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 181 67 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 181 67 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 67 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 67 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 67 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 179 67 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 179 67 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 67 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 67 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 67 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 177 67 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 177 67 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 67 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 67 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 67 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 175 67 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 175 67 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 174 67 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 174 67 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 28 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 28 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 27 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 27 67 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 26 67 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 26 67 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 26 67 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 25 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 25 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 24 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 24 67 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 198 67 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 197 67 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 197 67 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 67 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 67 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 196 67 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 195 67 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 195 67 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 67 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 67 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 194 67 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 193 67 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 193 67 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 67 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 67 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 192 67 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 191 67 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 191 67 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 67 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 67 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 190 67 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 189 67 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 189 67 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 67 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 67 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 188 67 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 187 67 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 187 67 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 67 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 67 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 186 67 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 185 67 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 185 67 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 67 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 67 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 184 67 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 183 67 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 183 67 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 67 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 67 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 182 67 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 181 67 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 181 67 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 67 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 67 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 180 67 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 179 67 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 179 67 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 67 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 67 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 178 67 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 177 67 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 177 67 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 67 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 67 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 176 67 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 175 67 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 175 67 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 174 67 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 67 174 67 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 28 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 28 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 27 67 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 27 67 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 26 67 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 26 67 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 26 67 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 25 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 25 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 24 67 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 24 67 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 198 66 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 197 66 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 197 66 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 196 66 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 196 66 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 196 66 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 195 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 195 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 194 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 194 66 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 194 66 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 193 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 193 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 192 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 192 66 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 192 66 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 191 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 191 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 190 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 190 66 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 190 66 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 189 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 189 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 188 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 188 66 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 188 66 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 187 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 187 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 186 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 186 66 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 186 66 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 185 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 185 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 184 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 184 66 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 184 66 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 183 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 183 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 182 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 182 66 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 182 66 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 181 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 181 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 180 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 180 66 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 180 66 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 179 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 179 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 178 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 178 66 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 178 66 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 177 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 177 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 176 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 176 66 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 176 66 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 175 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 175 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 174 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 174 66 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 28 66 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 28 66 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 27 66 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 27 66 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 26 66 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 26 66 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 26 66 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 25 66 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 25 66 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 24 66 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 24 66 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 198 66 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 197 66 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 197 66 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 196 66 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 196 66 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 196 66 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 195 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 195 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 194 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 194 66 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 194 66 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 193 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 193 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 192 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 192 66 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 192 66 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 191 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 191 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 190 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 190 66 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 190 66 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 189 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 189 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 188 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 188 66 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 188 66 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 187 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 187 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 186 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 186 66 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 186 66 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 185 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 185 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 184 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 184 66 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 184 66 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 183 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 183 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 182 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 182 66 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 182 66 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 181 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 181 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 180 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 180 66 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 180 66 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 179 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 179 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 178 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 178 66 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 178 66 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 177 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 177 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 176 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 176 66 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 176 66 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 175 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 175 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 174 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 66 174 66 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 28 66 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 28 66 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 27 66 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 27 66 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 66 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 66 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 66 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 25 66 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 25 66 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 24 66 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 24 66 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 198 66 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 197 66 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 197 66 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 66 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 66 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 66 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 195 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 195 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 66 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 66 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 66 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 193 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 193 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 66 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 66 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 66 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 191 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 191 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 66 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 66 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 66 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 189 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 189 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 66 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 66 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 66 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 187 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 187 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 66 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 66 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 66 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 185 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 185 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 66 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 66 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 66 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 183 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 183 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 66 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 66 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 66 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 181 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 181 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 66 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 66 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 66 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 179 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 179 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 66 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 66 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 66 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 177 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 177 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 66 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 66 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 66 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 175 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 175 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 174 66 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 174 66 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 28 65 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 28 65 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 27 65 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 27 65 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 65 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 65 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 65 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 25 65 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 25 65 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 24 65 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 24 65 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 198 65 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 197 65 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 197 65 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 65 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 65 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 65 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 195 65 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 195 65 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 65 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 65 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 65 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 193 65 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 193 65 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 65 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 65 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 65 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 191 65 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 191 65 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 65 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 65 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 65 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 189 65 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 189 65 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 65 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 65 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 65 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 187 65 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 187 65 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 65 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 65 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 65 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 185 65 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 185 65 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 65 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 65 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 65 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 183 65 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 183 65 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 65 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 65 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 65 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 181 65 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 181 65 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 65 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 65 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 65 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 179 65 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 179 65 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 65 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 65 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 65 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 177 65 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 177 65 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 65 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 65 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 65 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 175 65 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 175 65 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 174 65 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 174 65 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 28 65 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 28 65 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 27 65 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 27 65 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 65 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 65 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 26 65 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 25 65 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 25 65 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 24 65 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 24 65 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 198 65 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 197 65 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 197 65 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 65 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 65 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 196 65 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 195 65 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 195 65 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 65 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 65 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 194 65 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 193 65 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 193 65 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 65 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 65 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 192 65 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 191 65 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 191 65 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 65 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 65 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 190 65 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 189 65 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 189 65 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 65 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 65 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 188 65 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 187 65 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 187 65 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 65 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 65 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 186 65 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 185 65 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 185 65 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 65 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 65 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 184 65 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 183 65 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 183 65 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 65 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 65 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 182 65 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 181 65 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 181 65 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 65 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 65 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 180 65 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 179 65 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 179 65 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 65 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 65 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 178 65 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 177 65 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 177 65 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 65 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 65 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 176 65 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 175 65 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 175 65 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 174 65 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 65 174 65 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 28 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 28 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 27 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 27 64 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 26 64 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 26 64 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 26 64 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 25 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 25 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 24 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 24 64 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 198 64 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 197 64 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 197 64 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 196 64 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 196 64 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 196 64 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 195 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 195 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 194 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 194 64 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 194 64 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 193 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 193 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 192 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 192 64 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 192 64 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 191 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 191 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 190 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 190 64 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 190 64 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 189 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 189 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 188 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 188 64 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 188 64 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 187 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 187 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 186 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 186 64 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 186 64 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 185 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 185 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 184 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 184 64 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 184 64 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 183 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 183 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 182 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 182 64 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 182 64 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 181 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 181 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 180 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 180 64 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 180 64 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 179 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 179 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 178 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 178 64 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 178 64 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 177 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 177 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 176 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 176 64 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 176 64 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 175 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 175 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 174 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 174 64 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 28 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 28 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 27 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 27 64 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 26 64 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 26 64 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 26 64 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 25 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 25 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 24 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 24 64 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 198 64 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 197 64 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 197 64 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 196 64 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 196 64 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 196 64 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 195 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 195 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 194 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 194 64 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 194 64 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 193 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 193 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 192 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 192 64 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 192 64 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 191 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 191 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 190 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 190 64 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 190 64 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 189 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 189 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 188 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 188 64 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 188 64 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 187 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 187 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 186 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 186 64 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 186 64 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 185 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 185 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 184 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 184 64 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 184 64 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 183 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 183 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 182 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 182 64 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 182 64 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 181 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 181 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 180 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 180 64 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 180 64 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 179 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 179 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 178 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 178 64 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 178 64 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 177 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 177 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 176 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 176 64 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 176 64 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 175 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 175 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 174 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 64 174 64 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 28 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 28 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 27 64 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 27 64 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 64 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 64 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 64 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 25 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 25 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 24 64 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 24 64 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 198 64 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 197 64 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 197 64 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 64 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 64 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 64 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 195 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 195 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 64 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 64 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 64 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 193 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 193 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 64 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 64 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 64 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 191 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 191 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 64 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 64 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 64 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 189 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 189 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 64 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 64 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 64 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 187 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 187 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 64 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 64 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 64 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 185 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 185 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 64 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 64 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 64 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 183 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 183 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 64 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 64 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 64 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 181 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 181 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 64 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 64 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 64 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 179 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 179 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 64 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 64 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 64 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 177 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 177 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 64 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 64 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 64 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 175 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 175 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 174 64 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 174 64 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 28 63 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 28 63 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 27 63 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 27 63 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 63 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 63 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 63 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 25 63 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 25 63 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 24 63 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 24 63 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 198 63 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 197 63 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 197 63 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 63 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 63 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 63 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 195 63 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 195 63 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 63 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 63 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 63 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 193 63 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 193 63 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 63 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 63 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 63 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 191 63 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 191 63 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 63 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 63 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 63 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 189 63 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 189 63 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 63 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 63 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 63 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 187 63 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 187 63 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 63 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 63 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 63 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 185 63 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 185 63 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 63 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 63 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 63 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 183 63 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 183 63 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 63 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 63 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 63 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 181 63 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 181 63 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 63 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 63 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 63 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 179 63 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 179 63 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 63 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 63 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 63 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 177 63 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 177 63 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 63 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 63 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 63 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 175 63 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 175 63 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 174 63 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 174 63 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 28 63 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 28 63 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 27 63 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 27 63 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 63 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 63 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 26 63 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 25 63 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 25 63 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 24 63 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 24 63 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 198 63 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 197 63 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 197 63 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 63 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 63 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 196 63 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 195 63 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 195 63 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 63 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 63 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 194 63 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 193 63 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 193 63 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 63 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 63 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 192 63 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 191 63 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 191 63 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 63 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 63 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 190 63 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 189 63 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 189 63 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 63 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 63 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 188 63 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 187 63 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 187 63 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 63 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 63 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 186 63 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 185 63 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 185 63 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 63 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 63 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 184 63 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 183 63 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 183 63 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 63 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 63 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 182 63 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 181 63 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 181 63 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 63 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 63 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 180 63 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 179 63 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 179 63 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 63 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 63 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 178 63 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 177 63 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 177 63 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 63 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 63 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 176 63 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 175 63 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 175 63 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 174 63 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 63 174 63 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 28 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 28 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 27 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 27 62 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 26 62 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 26 62 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 26 62 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 25 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 25 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 24 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 24 62 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 198 62 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 197 62 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 197 62 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 196 62 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 196 62 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 196 62 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 195 62 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 195 62 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 194 62 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 194 62 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 194 62 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 193 62 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 193 62 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 192 62 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 192 62 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 192 62 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 191 62 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 191 62 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 190 62 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 190 62 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 190 62 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 189 62 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 189 62 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 188 62 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 188 62 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 188 62 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 187 62 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 187 62 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 186 62 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 186 62 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 186 62 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 185 62 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 185 62 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 184 62 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 184 62 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 184 62 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 183 62 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 183 62 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 182 62 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 182 62 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 182 62 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 181 62 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 181 62 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 180 62 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 180 62 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 180 62 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 179 62 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 179 62 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 178 62 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 178 62 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 178 62 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 177 62 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 177 62 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 176 62 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 176 62 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 176 62 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 175 62 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 175 62 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 174 62 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 174 62 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 28 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 28 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 27 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 27 62 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 26 62 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 26 62 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 26 62 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 25 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 25 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 24 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 62 24 62 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 28 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 28 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 27 62 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 27 62 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 62 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 62 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 62 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 25 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 25 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 24 62 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 24 62 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 28 61 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 28 61 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 27 61 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 27 61 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 61 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 61 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 61 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 25 61 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 25 61 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 24 61 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 24 61 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 28 61 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 28 61 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 27 61 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 27 61 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 61 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 61 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 26 61 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 25 61 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 25 61 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 24 61 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 61 24 61 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 28 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 28 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 27 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 27 60 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 26 60 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 26 60 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 26 60 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 25 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 25 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 24 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 24 60 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 28 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 28 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 27 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 27 60 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 26 60 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 26 60 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 26 60 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 25 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 25 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 24 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 60 24 60 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 28 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 28 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 27 60 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 27 60 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 60 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 60 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 60 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 25 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 25 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 24 60 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 24 60 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 28 59 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 28 59 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 27 59 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 27 59 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 59 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 59 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 59 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 25 59 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 25 59 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 24 59 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 24 59 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 28 59 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 28 59 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 27 59 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 27 59 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 59 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 59 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 26 59 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 25 59 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 25 59 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 24 59 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 59 24 59 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 28 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 28 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 27 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 27 58 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 26 58 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 26 58 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 26 58 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 25 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 25 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 24 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 24 58 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 28 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 28 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 27 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 27 58 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 26 58 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 26 58 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 26 58 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 25 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 25 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 24 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 58 24 58 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 28 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 28 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 27 58 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 27 58 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 58 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 58 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 58 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 25 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 25 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 24 58 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 24 58 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 28 57 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 28 57 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 27 57 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 27 57 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 57 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 57 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 57 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 25 57 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 25 57 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 24 57 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 24 57 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 28 57 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 28 57 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 27 57 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 27 57 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 57 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 57 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 26 57 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 25 57 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 25 57 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 24 57 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 57 24 57 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 28 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 28 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 27 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 27 56 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 26 56 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 26 56 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 26 56 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 25 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 25 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 24 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 24 56 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 28 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 28 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 27 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 27 56 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 26 56 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 26 56 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 26 56 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 25 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 25 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 24 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 56 24 56 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 28 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 28 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 27 56 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 27 56 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 56 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 56 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 56 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 25 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 25 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 24 56 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 24 56 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 28 55 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 28 55 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 27 55 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 27 55 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 55 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 55 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 55 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 25 55 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 25 55 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 24 55 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 24 55 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 28 55 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 28 55 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 27 55 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 27 55 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 55 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 55 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 26 55 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 25 55 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 25 55 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 24 55 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 55 24 55 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 28 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 28 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 27 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 27 54 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 26 54 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 26 54 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 26 54 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 25 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 25 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 24 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 24 54 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 28 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 28 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 27 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 27 54 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 26 54 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 26 54 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 26 54 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 25 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 25 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 24 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 54 24 54 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 28 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 28 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 27 54 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 27 54 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 26 54 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 26 54 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 26 54 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 25 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 25 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 24 54 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 24 54 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 28 53 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 28 53 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 27 53 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 27 53 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 26 53 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 26 53 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 26 53 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 25 53 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 25 53 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 24 53 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 53 24 53 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 28 53 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 28 53 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 27 53 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 27 53 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 53 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 53 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 53 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 25 53 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 25 53 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 24 53 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 24 53 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 28 52 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 28 52 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 27 52 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 27 52 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 52 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 52 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 52 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 25 52 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 25 52 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 24 52 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 24 52 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 28 52 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 28 52 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 27 52 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 27 52 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 52 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 52 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 26 52 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 25 52 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 25 52 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 24 52 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 52 24 52 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 28 51 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 28 51 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 27 51 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 27 51 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 26 51 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 26 51 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 26 51 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 25 51 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 25 51 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 24 51 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 24 51 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 28 51 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 28 51 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 27 51 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 27 51 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 26 51 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 26 51 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 26 51 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 25 51 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 25 51 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 24 51 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 51 24 51 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 28 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 28 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 27 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 27 24 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 26 24 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 26 24 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 26 24 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 25 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 25 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 24 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 24 24 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 28 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 28 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 27 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 27 24 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 26 24 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 26 24 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 26 24 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 25 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 25 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 24 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 24 24 24 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 28 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 28 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 27 24 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 27 24 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 26 24 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 26 24 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 26 24 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 25 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 25 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 24 24 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 24 24 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 28 23 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 28 23 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 27 23 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 27 23 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 26 23 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 26 23 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 26 23 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 25 23 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 25 23 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 24 23 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 23 24 23 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 28 23 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 28 23 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 27 23 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 27 23 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 23 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 23 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 23 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 25 23 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 25 23 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 24 23 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 24 23 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 28 22 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 28 22 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 27 22 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 27 22 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 22 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 22 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 22 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 25 22 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 25 22 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 24 22 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 24 22 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 28 22 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 28 22 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 27 22 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 27 22 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 22 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 22 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 26 22 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 25 22 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 25 22 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 24 22 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 22 24 22 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 28 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 28 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 27 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 27 21 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 26 21 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 26 21 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 26 21 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 25 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 25 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 24 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 24 21 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 28 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 28 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 27 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 27 21 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 26 21 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 26 21 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 26 21 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 25 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 25 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 24 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 21 24 21 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 28 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 28 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 27 21 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 27 21 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 21 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 21 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 21 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 25 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 25 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 24 21 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 24 21 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 28 20 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 28 20 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 27 20 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 27 20 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 20 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 20 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 20 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 25 20 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 25 20 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 24 20 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 24 20 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 28 20 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 28 20 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 27 20 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 27 20 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 20 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 20 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 26 20 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 25 20 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 25 20 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 24 20 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 20 24 20 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 28 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 28 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 27 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 27 19 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 26 19 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 26 19 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 26 19 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 25 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 25 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 24 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 24 19 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 28 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 28 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 27 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 27 19 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 26 19 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 26 19 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 26 19 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 25 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 25 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 24 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 19 24 19 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 28 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 28 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 27 19 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 27 19 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 19 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 19 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 19 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 25 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 25 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 24 19 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 24 19 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 28 18 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 28 18 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 27 18 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 27 18 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 18 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 18 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 18 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 25 18 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 25 18 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 24 18 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 24 18 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 28 18 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 28 18 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 27 18 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 27 18 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 18 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 18 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 26 18 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 25 18 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 25 18 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 24 18 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 18 24 18 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 28 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 28 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 27 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 27 17 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 26 17 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 26 17 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 26 17 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 25 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 25 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 24 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 24 17 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 28 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 28 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 27 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 27 17 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 26 17 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 26 17 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 26 17 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 25 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 25 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 24 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 17 24 17 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 28 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 28 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 27 17 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 27 17 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 17 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 17 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 17 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 25 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 25 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 24 17 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 24 17 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 28 16 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 28 16 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 27 16 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 27 16 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 16 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 16 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 16 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 25 16 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 25 16 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 24 16 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 24 16 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 28 16 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 28 16 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 27 16 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 27 16 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 16 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 16 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 26 16 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 25 16 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 25 16 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 24 16 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 16 24 16 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 28 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 28 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 27 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 27 15 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 26 15 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 26 15 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 26 15 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 25 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 25 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 24 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 24 15 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 28 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 28 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 27 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 27 15 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 26 15 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 26 15 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 26 15 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 25 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 25 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 24 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 15 24 15 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 28 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 28 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 27 15 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 27 15 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 15 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 15 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 15 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 25 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 25 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 24 15 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 24 15 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 28 14 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 28 14 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 27 14 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 27 14 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 14 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 14 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 14 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 25 14 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 25 14 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 24 14 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 24 14 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 28 14 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 28 14 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 27 14 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 27 14 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 14 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 14 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 26 14 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 25 14 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 25 14 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 24 14 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 14 24 14 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 28 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 28 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 27 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 27 13 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 26 13 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 26 13 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 26 13 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 25 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 25 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 24 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 24 13 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 28 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 28 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 27 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 27 13 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 26 13 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 26 13 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 26 13 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 25 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 25 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 24 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 24 13 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 198 13 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 197 13 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 197 13 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 196 13 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 196 13 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 196 13 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 195 13 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 195 13 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 194 13 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 194 13 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 194 13 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 193 13 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 193 13 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 192 13 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 192 13 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 192 13 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 191 13 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 191 13 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 190 13 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 190 13 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 190 13 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 189 13 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 189 13 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 188 13 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 188 13 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 188 13 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 187 13 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 187 13 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 186 13 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 186 13 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 186 13 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 185 13 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 185 13 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 184 13 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 184 13 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 184 13 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 183 13 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 183 13 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 182 13 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 182 13 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 182 13 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 181 13 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 181 13 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 180 13 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 180 13 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 180 13 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 179 13 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 179 13 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 178 13 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 178 13 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 178 13 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 177 13 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 177 13 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 176 13 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 176 13 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 176 13 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 175 13 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 175 13 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 174 13 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 13 174 13 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 28 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 28 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 27 13 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 27 13 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 13 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 13 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 13 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 25 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 25 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 24 13 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 24 13 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 198 12 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 197 12 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 197 12 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 196 12 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 196 12 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 196 12 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 195 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 195 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 194 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 194 12 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 194 12 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 193 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 193 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 192 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 192 12 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 192 12 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 191 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 191 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 190 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 190 12 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 190 12 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 189 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 189 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 188 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 188 12 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 188 12 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 187 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 187 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 186 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 186 12 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 186 12 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 185 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 185 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 184 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 184 12 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 184 12 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 183 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 183 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 182 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 182 12 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 182 12 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 181 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 181 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 180 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 180 12 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 180 12 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 179 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 179 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 178 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 178 12 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 178 12 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 177 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 177 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 176 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 176 12 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 176 12 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 175 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 175 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 174 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 174 12 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 28 12 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 28 12 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 27 12 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 27 12 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 12 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 12 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 12 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 25 12 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 25 12 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 24 12 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 24 12 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 198 12 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 197 12 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 197 12 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 196 12 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 196 12 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 196 12 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 195 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 195 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 194 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 194 12 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 194 12 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 193 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 193 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 192 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 192 12 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 192 12 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 191 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 191 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 190 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 190 12 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 190 12 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 189 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 189 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 188 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 188 12 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 188 12 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 187 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 187 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 186 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 186 12 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 186 12 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 185 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 185 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 184 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 184 12 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 184 12 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 183 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 183 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 182 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 182 12 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 182 12 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 181 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 181 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 180 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 180 12 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 180 12 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 179 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 179 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 178 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 178 12 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 178 12 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 177 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 177 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 176 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 176 12 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 176 12 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 175 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 175 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 174 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 174 12 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 28 12 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 28 12 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 27 12 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 27 12 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 12 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 12 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 26 12 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 25 12 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 25 12 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 24 12 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 12 24 12 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 198 12 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 197 12 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 197 12 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 12 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 12 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 12 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 195 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 195 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 12 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 12 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 12 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 193 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 193 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 12 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 12 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 12 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 191 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 191 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 12 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 12 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 12 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 189 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 189 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 12 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 12 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 12 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 187 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 187 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 12 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 12 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 12 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 185 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 185 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 12 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 12 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 12 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 183 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 183 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 12 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 12 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 12 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 181 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 181 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 12 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 12 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 12 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 179 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 179 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 12 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 12 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 12 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 177 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 177 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 12 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 12 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 12 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 175 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 175 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 174 12 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 174 12 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 28 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 28 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 27 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 27 11 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 26 11 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 26 11 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 26 11 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 25 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 25 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 24 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 24 11 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 198 11 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 197 11 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 197 11 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 11 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 11 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 11 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 195 11 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 195 11 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 11 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 11 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 11 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 193 11 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 193 11 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 11 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 11 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 11 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 191 11 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 191 11 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 11 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 11 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 11 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 189 11 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 189 11 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 11 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 11 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 11 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 187 11 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 187 11 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 11 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 11 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 11 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 185 11 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 185 11 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 11 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 11 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 11 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 183 11 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 183 11 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 11 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 11 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 11 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 181 11 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 181 11 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 11 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 11 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 11 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 179 11 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 179 11 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 11 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 11 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 11 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 177 11 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 177 11 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 11 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 11 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 11 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 175 11 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 175 11 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 174 11 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 174 11 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 28 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 28 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 27 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 27 11 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 26 11 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 26 11 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 26 11 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 25 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 25 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 24 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 24 11 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 198 11 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 197 11 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 197 11 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 11 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 11 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 196 11 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 195 11 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 195 11 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 11 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 11 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 194 11 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 193 11 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 193 11 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 11 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 11 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 192 11 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 191 11 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 191 11 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 11 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 11 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 190 11 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 189 11 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 189 11 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 11 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 11 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 188 11 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 187 11 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 187 11 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 11 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 11 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 186 11 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 185 11 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 185 11 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 11 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 11 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 184 11 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 183 11 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 183 11 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 11 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 11 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 182 11 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 181 11 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 181 11 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 11 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 11 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 180 11 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 179 11 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 179 11 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 11 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 11 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 178 11 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 177 11 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 177 11 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 11 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 11 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 176 11 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 175 11 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 175 11 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 174 11 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 11 174 11 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 28 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 28 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 27 11 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 27 11 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 11 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 11 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 11 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 25 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 25 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 24 11 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 24 11 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 198 10 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 197 10 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 197 10 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 196 10 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 196 10 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 196 10 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 195 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 195 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 194 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 194 10 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 194 10 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 193 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 193 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 192 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 192 10 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 192 10 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 191 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 191 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 190 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 190 10 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 190 10 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 189 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 189 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 188 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 188 10 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 188 10 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 187 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 187 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 186 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 186 10 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 186 10 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 185 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 185 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 184 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 184 10 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 184 10 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 183 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 183 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 182 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 182 10 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 182 10 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 181 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 181 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 180 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 180 10 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 180 10 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 179 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 179 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 178 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 178 10 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 178 10 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 177 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 177 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 176 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 176 10 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 176 10 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 175 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 175 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 174 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 174 10 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 28 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 28 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 27 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 27 10 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 10 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 10 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 10 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 25 10 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 25 10 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 24 10 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 24 10 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 198 10 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 197 10 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 197 10 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 196 10 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 196 10 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 196 10 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 195 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 195 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 194 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 194 10 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 194 10 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 193 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 193 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 192 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 192 10 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 192 10 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 191 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 191 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 190 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 190 10 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 190 10 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 189 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 189 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 188 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 188 10 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 188 10 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 187 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 187 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 186 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 186 10 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 186 10 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 185 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 185 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 184 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 184 10 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 184 10 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 183 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 183 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 182 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 182 10 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 182 10 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 181 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 181 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 180 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 180 10 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 180 10 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 179 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 179 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 178 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 178 10 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 178 10 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 177 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 177 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 176 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 176 10 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 176 10 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 175 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 175 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 174 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 174 10 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 28 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 28 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 27 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 27 10 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 10 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 10 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 26 10 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 25 10 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 25 10 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 24 10 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 10 24 10 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 198 10 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 197 10 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 197 10 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 10 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 10 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 10 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 195 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 195 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 10 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 10 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 10 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 193 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 193 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 10 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 10 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 10 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 191 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 191 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 10 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 10 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 10 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 189 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 189 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 10 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 10 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 10 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 187 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 187 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 10 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 10 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 10 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 185 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 185 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 10 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 10 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 10 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 183 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 183 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 10 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 10 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 10 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 181 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 181 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 10 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 10 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 10 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 179 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 179 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 10 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 10 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 10 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 177 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 177 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 10 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 10 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 10 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 175 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 175 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 174 10 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 174 10 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 28 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 28 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 27 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 27 9 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 26 9 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 26 9 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 26 9 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 25 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 25 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 24 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 24 9 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 198 9 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 197 9 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 197 9 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 9 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 9 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 9 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 195 9 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 195 9 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 9 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 9 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 9 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 193 9 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 193 9 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 9 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 9 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 9 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 191 9 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 191 9 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 9 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 9 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 9 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 189 9 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 189 9 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 9 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 9 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 9 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 187 9 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 187 9 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 9 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 9 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 9 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 185 9 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 185 9 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 9 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 9 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 9 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 183 9 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 183 9 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 9 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 9 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 9 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 181 9 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 181 9 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 9 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 9 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 9 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 179 9 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 179 9 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 9 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 9 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 9 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 177 9 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 177 9 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 9 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 9 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 9 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 175 9 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 175 9 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 174 9 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 174 9 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 28 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 28 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 27 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 27 9 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 26 9 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 26 9 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 26 9 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 25 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 25 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 24 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 24 9 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 198 9 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 197 9 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 197 9 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 9 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 9 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 196 9 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 195 9 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 195 9 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 9 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 9 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 194 9 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 193 9 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 193 9 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 9 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 9 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 192 9 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 191 9 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 191 9 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 9 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 9 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 190 9 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 189 9 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 189 9 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 9 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 9 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 188 9 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 187 9 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 187 9 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 9 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 9 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 186 9 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 185 9 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 185 9 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 9 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 9 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 184 9 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 183 9 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 183 9 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 9 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 9 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 182 9 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 181 9 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 181 9 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 9 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 9 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 180 9 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 179 9 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 179 9 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 9 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 9 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 178 9 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 177 9 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 177 9 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 9 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 9 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 176 9 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 175 9 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 175 9 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 174 9 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 9 174 9 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 28 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 28 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 27 9 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 27 9 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 9 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 9 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 9 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 25 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 25 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 24 9 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 24 9 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 198 8 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 197 8 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 197 8 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 196 8 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 196 8 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 196 8 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 195 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 195 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 194 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 194 8 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 194 8 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 193 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 193 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 192 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 192 8 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 192 8 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 191 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 191 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 190 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 190 8 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 190 8 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 189 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 189 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 188 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 188 8 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 188 8 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 187 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 187 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 186 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 186 8 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 186 8 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 185 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 185 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 184 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 184 8 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 184 8 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 183 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 183 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 182 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 182 8 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 182 8 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 181 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 181 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 180 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 180 8 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 180 8 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 179 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 179 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 178 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 178 8 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 178 8 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 177 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 177 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 176 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 176 8 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 176 8 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 175 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 175 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 174 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 174 8 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 28 8 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 28 8 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 27 8 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 27 8 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 8 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 8 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 8 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 25 8 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 25 8 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 24 8 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 24 8 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 198 8 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 197 8 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 197 8 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 196 8 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 196 8 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 196 8 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 195 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 195 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 194 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 194 8 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 194 8 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 193 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 193 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 192 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 192 8 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 192 8 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 191 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 191 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 190 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 190 8 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 190 8 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 189 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 189 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 188 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 188 8 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 188 8 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 187 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 187 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 186 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 186 8 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 186 8 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 185 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 185 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 184 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 184 8 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 184 8 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 183 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 183 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 182 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 182 8 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 182 8 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 181 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 181 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 180 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 180 8 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 180 8 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 179 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 179 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 178 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 178 8 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 178 8 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 177 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 177 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 176 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 176 8 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 176 8 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 175 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 175 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 174 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 174 8 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 28 8 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 28 8 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 27 8 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 27 8 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 8 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 8 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 26 8 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 25 8 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 25 8 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 24 8 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 8 24 8 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 198 8 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 197 8 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 197 8 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 8 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 8 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 8 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 195 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 195 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 8 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 8 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 8 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 193 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 193 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 8 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 8 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 8 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 191 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 191 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 8 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 8 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 8 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 189 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 189 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 8 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 8 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 8 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 187 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 187 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 8 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 8 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 8 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 185 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 185 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 8 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 8 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 8 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 183 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 183 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 8 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 8 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 8 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 181 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 181 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 8 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 8 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 8 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 179 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 179 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 8 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 8 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 8 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 177 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 177 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 8 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 8 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 8 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 175 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 175 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 174 8 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 174 8 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 28 7 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 28 7 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 27 7 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 27 7 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 26 7 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 26 7 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 26 7 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 25 7 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 25 7 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 24 7 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 24 7 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 198 7 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 197 7 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 197 7 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 7 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 7 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 7 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 195 7 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 195 7 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 7 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 7 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 7 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 193 7 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 193 7 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 7 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 7 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 7 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 191 7 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 191 7 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 7 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 7 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 7 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 189 7 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 189 7 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 7 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 7 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 7 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 187 7 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 187 7 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 7 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 7 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 7 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 185 7 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 185 7 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 7 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 7 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 7 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 183 7 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 183 7 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 7 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 7 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 7 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 181 7 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 181 7 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 7 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 7 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 7 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 179 7 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 179 7 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 7 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 7 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 7 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 177 7 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 177 7 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 7 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 7 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 7 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 175 7 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 175 7 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 174 7 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 174 7 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 28 7 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 28 7 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 27 7 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 27 7 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 26 7 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 26 7 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 26 7 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 25 7 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 25 7 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 24 7 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 24 7 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 198 7 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 197 7 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 197 7 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 7 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 7 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 196 7 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 195 7 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 195 7 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 7 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 7 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 194 7 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 193 7 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 193 7 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 7 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 7 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 192 7 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 191 7 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 191 7 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 7 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 7 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 190 7 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 189 7 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 189 7 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 7 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 7 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 188 7 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 187 7 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 187 7 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 7 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 7 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 186 7 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 185 7 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 185 7 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 7 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 7 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 184 7 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 183 7 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 183 7 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 7 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 7 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 182 7 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 181 7 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 181 7 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 7 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 7 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 180 7 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 179 7 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 179 7 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 7 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 7 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 178 7 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 177 7 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 177 7 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 7 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 7 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 176 7 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 175 7 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 175 7 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 174 7 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 7 174 7 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 28 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 28 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 27 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 27 6 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 26 6 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 26 6 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 26 6 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 25 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 25 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 24 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 24 6 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 198 6 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 197 6 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 197 6 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 196 6 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 196 6 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 196 6 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 195 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 195 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 194 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 194 6 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 194 6 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 193 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 193 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 192 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 192 6 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 192 6 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 191 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 191 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 190 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 190 6 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 190 6 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 189 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 189 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 188 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 188 6 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 188 6 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 187 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 187 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 186 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 186 6 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 186 6 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 185 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 185 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 184 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 184 6 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 184 6 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 183 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 183 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 182 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 182 6 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 182 6 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 181 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 181 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 180 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 180 6 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 180 6 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 179 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 179 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 178 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 178 6 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 178 6 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 177 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 177 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 176 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 176 6 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 176 6 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 175 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 175 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 174 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 174 6 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 28 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 28 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 27 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 27 6 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 26 6 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 26 6 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 26 6 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 25 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 25 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 24 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 24 6 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 198 6 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 197 6 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 197 6 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 196 6 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 196 6 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 196 6 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 195 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 195 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 194 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 194 6 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 194 6 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 193 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 193 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 192 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 192 6 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 192 6 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 191 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 191 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 190 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 190 6 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 190 6 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 189 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 189 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 188 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 188 6 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 188 6 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 187 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 187 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 186 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 186 6 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 186 6 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 185 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 185 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 184 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 184 6 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 184 6 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 183 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 183 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 182 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 182 6 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 182 6 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 181 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 181 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 180 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 180 6 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 180 6 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 179 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 179 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 178 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 178 6 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 178 6 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 177 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 177 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 176 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 176 6 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 176 6 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 175 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 175 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 174 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 6 174 6 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 28 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 28 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 27 6 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 27 6 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 6 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 6 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 6 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 25 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 25 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 24 6 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 24 6 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 198 6 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 197 6 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 197 6 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 6 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 6 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 6 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 195 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 195 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 6 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 6 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 6 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 193 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 193 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 6 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 6 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 6 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 191 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 191 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 6 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 6 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 6 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 189 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 189 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 6 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 6 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 6 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 187 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 187 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 6 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 6 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 6 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 185 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 185 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 6 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 6 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 6 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 183 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 183 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 6 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 6 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 6 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 181 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 181 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 6 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 6 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 6 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 179 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 179 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 6 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 6 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 6 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 177 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 177 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 6 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 6 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 6 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 175 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 175 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 174 6 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 174 6 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 28 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 28 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 27 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 27 5 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 5 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 5 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 5 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 25 5 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 25 5 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 24 5 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 24 5 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 198 5 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 197 5 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 197 5 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 5 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 5 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 5 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 195 5 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 195 5 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 5 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 5 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 5 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 193 5 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 193 5 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 5 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 5 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 5 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 191 5 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 191 5 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 5 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 5 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 5 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 189 5 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 189 5 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 5 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 5 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 5 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 187 5 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 187 5 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 5 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 5 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 5 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 185 5 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 185 5 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 5 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 5 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 5 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 183 5 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 183 5 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 5 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 5 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 5 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 181 5 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 181 5 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 5 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 5 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 5 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 179 5 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 179 5 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 5 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 5 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 5 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 177 5 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 177 5 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 5 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 5 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 5 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 175 5 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 175 5 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 174 5 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 174 5 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 28 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 28 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 27 5 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 27 5 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 5 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 5 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 26 5 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 25 5 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 25 5 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 24 5 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 24 5 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 198 5 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 197 5 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 197 5 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 5 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 5 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 196 5 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 195 5 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 195 5 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 5 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 5 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 194 5 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 193 5 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 193 5 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 5 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 5 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 192 5 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 191 5 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 191 5 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 5 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 5 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 190 5 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 189 5 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 189 5 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 5 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 5 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 188 5 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 187 5 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 187 5 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 5 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 5 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 186 5 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 185 5 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 185 5 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 5 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 5 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 184 5 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 183 5 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 183 5 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 5 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 5 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 182 5 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 181 5 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 181 5 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 5 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 5 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 180 5 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 179 5 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 179 5 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 5 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 5 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 178 5 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 177 5 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 177 5 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 5 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 5 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 176 5 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 175 5 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 175 5 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 174 5 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 5 174 5 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 28 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 28 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 27 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 27 4 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 26 4 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 26 4 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 26 4 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 25 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 25 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 24 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 24 4 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 198 4 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 197 4 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 197 4 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 196 4 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 196 4 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 196 4 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 195 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 195 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 194 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 194 4 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 194 4 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 193 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 193 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 192 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 192 4 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 192 4 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 191 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 191 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 190 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 190 4 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 190 4 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 189 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 189 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 188 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 188 4 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 188 4 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 187 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 187 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 186 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 186 4 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 186 4 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 185 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 185 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 184 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 184 4 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 184 4 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 183 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 183 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 182 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 182 4 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 182 4 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 181 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 181 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 180 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 180 4 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 180 4 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 179 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 179 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 178 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 178 4 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 178 4 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 177 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 177 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 176 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 176 4 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 176 4 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 175 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 175 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 174 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 174 4 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 28 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 28 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 27 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 27 4 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 26 4 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 26 4 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 26 4 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 25 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 25 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 24 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 24 4 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 198 4 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 197 4 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 197 4 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 196 4 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 196 4 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 196 4 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 195 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 195 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 194 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 194 4 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 194 4 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 193 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 193 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 192 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 192 4 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 192 4 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 191 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 191 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 190 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 190 4 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 190 4 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 189 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 189 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 188 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 188 4 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 188 4 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 187 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 187 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 186 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 186 4 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 186 4 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 185 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 185 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 184 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 184 4 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 184 4 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 183 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 183 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 182 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 182 4 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 182 4 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 181 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 181 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 180 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 180 4 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 180 4 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 179 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 179 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 178 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 178 4 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 178 4 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 177 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 177 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 176 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 176 4 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 176 4 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 175 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 175 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 174 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 4 174 4 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 28 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 28 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 27 4 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 27 4 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 4 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 4 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 4 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 25 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 25 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 24 4 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 24 4 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 198 4 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 197 4 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 197 4 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 4 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 4 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 4 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 195 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 195 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 4 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 4 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 4 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 193 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 193 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 4 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 4 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 4 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 191 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 191 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 4 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 4 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 4 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 189 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 189 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 4 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 4 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 4 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 187 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 187 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 4 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 4 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 4 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 185 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 185 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 4 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 4 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 4 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 183 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 183 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 4 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 4 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 4 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 181 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 181 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 4 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 4 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 4 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 179 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 179 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 4 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 4 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 4 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 177 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 177 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 4 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 4 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 4 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 175 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 175 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 174 4 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 174 4 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 28 3 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 28 3 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 27 3 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 27 3 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 3 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 3 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 3 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 25 3 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 25 3 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 24 3 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 24 3 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 198 3 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 197 3 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 197 3 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 3 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 3 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 3 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 195 3 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 195 3 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 3 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 3 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 3 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 193 3 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 193 3 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 3 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 3 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 3 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 191 3 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 191 3 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 3 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 3 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 3 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 189 3 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 189 3 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 3 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 3 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 3 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 187 3 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 187 3 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 3 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 3 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 3 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 185 3 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 185 3 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 3 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 3 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 3 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 183 3 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 183 3 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 3 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 3 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 3 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 181 3 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 181 3 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 3 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 3 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 3 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 179 3 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 179 3 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 3 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 3 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 3 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 177 3 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 177 3 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 3 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 3 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 3 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 175 3 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 175 3 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 174 3 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 174 3 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 28 3 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 28 3 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 27 3 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 27 3 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 3 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 3 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 26 3 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 25 3 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 25 3 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 24 3 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 24 3 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 198 3 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 197 3 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 197 3 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 3 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 3 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 196 3 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 195 3 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 195 3 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 3 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 3 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 194 3 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 193 3 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 193 3 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 3 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 3 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 192 3 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 191 3 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 191 3 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 3 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 3 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 190 3 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 189 3 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 189 3 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 3 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 3 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 188 3 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 187 3 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 187 3 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 3 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 3 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 186 3 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 185 3 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 185 3 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 3 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 3 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 184 3 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 183 3 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 183 3 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 3 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 3 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 182 3 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 181 3 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 181 3 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 3 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 3 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 180 3 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 179 3 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 179 3 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 3 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 3 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 178 3 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 177 3 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 177 3 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 3 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 3 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 176 3 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 175 3 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 175 3 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 174 3 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 3 174 3 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 28 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 28 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 27 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 27 2 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 26 2 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 26 2 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 26 2 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 25 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 25 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 24 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 24 2 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 198 2 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 197 2 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 197 2 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 196 2 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 196 2 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 196 2 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 195 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 195 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 194 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 194 2 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 194 2 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 193 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 193 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 192 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 192 2 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 192 2 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 191 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 191 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 190 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 190 2 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 190 2 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 189 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 189 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 188 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 188 2 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 188 2 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 187 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 187 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 186 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 186 2 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 186 2 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 185 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 185 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 184 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 184 2 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 184 2 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 183 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 183 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 182 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 182 2 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 182 2 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 181 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 181 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 180 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 180 2 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 180 2 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 179 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 179 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 178 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 178 2 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 178 2 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 177 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 177 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 176 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 176 2 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 176 2 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 175 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 175 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 174 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 174 2 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 28 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 28 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 27 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 27 2 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 26 2 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 26 2 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 26 2 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 25 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 25 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 24 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 24 2 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 198 2 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 197 2 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 197 2 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 196 2 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 196 2 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 196 2 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 195 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 195 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 194 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 194 2 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 194 2 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 193 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 193 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 192 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 192 2 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 192 2 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 191 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 191 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 190 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 190 2 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 190 2 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 189 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 189 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 188 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 188 2 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 188 2 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 187 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 187 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 186 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 186 2 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 186 2 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 185 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 185 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 184 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 184 2 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 184 2 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 183 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 183 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 182 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 182 2 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 182 2 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 181 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 181 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 180 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 180 2 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 180 2 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 179 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 179 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 178 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 178 2 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 178 2 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 177 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 177 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 176 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 176 2 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 176 2 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 175 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 175 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 174 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 2 174 2 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 198 2 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 197 2 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 197 2 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 2 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 2 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 2 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 195 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 195 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 2 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 2 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 2 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 193 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 193 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 2 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 2 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 2 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 191 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 191 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 2 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 2 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 2 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 189 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 189 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 2 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 2 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 2 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 187 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 187 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 2 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 2 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 2 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 185 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 185 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 2 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 2 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 2 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 183 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 183 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 2 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 2 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 2 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 181 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 181 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 2 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 2 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 2 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 179 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 179 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 2 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 2 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 2 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 177 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 177 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 2 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 2 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 2 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 175 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 175 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 174 2 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 174 2 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 28 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 28 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 27 2 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 27 2 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 2 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 2 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 2 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 25 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 25 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 24 2 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 24 2 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 198 1 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 197 1 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 197 1 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 1 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 1 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 1 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 195 1 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 195 1 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 1 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 1 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 1 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 193 1 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 193 1 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 1 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 1 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 1 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 191 1 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 191 1 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 1 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 1 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 1 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 189 1 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 189 1 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 1 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 1 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 1 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 187 1 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 187 1 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 1 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 1 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 1 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 185 1 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 185 1 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 1 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 1 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 1 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 183 1 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 183 1 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 1 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 1 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 1 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 181 1 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 181 1 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 1 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 1 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 1 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 179 1 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 179 1 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 1 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 1 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 1 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 177 1 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 177 1 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 1 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 1 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 1 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 175 1 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 175 1 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 174 1 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 174 1 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 28 1 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 28 1 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 27 1 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 27 1 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 1 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 1 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 1 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 25 1 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 25 1 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 24 1 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 24 1 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 198 1 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 197 1 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 197 1 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 1 197 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 1 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 196 1 196 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 195 1 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 195 1 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 1 195 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 1 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 194 1 194 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 193 1 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 193 1 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 1 193 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 1 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 192 1 192 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 191 1 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 191 1 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 1 191 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 1 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 190 1 190 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 189 1 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 189 1 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 1 189 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 1 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 188 1 188 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 187 1 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 187 1 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 1 187 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 1 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 186 1 186 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 185 1 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 185 1 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 1 185 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 1 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 184 1 184 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 183 1 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 183 1 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 1 183 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 1 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 182 1 182 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 181 1 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 181 1 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 1 181 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 1 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 180 1 180 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 179 1 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 179 1 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 1 179 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 1 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 178 1 178 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 177 1 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 177 1 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 1 177 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 1 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 176 1 176 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 175 1 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 175 1 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 174 1 175 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 174 1 174 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 28 1 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 28 1 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 27 1 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 27 1 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 1 27 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 1 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 26 1 26 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 25 1 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 25 1 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 24 1 25 6 VSSIO
port 10 nsew ground bidirectional
rlabel nfet_brown s 1 24 1 24 6 VSSIO
port 10 nsew ground bidirectional
rlabel 
 s 1 56 24 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel 
 s 51 56 74 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 56 24 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 51 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 60 74 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 60 74 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 60 74 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 59 74 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 59 74 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 58 74 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 58 74 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 58 74 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 57 74 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 57 74 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 56 74 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 60 74 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 60 74 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 60 74 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 59 74 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 59 74 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 58 74 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 58 74 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 58 74 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 57 74 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 57 74 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 74 56 74 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 60 73 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 60 73 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 60 73 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 59 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 59 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 58 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 58 73 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 58 73 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 57 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 57 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 56 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 60 73 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 60 73 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 60 73 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 59 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 59 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 58 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 58 73 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 58 73 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 57 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 57 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 73 56 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 73 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 73 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 73 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 59 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 59 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 73 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 73 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 73 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 57 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 57 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 56 73 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 72 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 72 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 72 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 59 72 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 59 72 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 72 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 72 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 72 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 57 72 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 57 72 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 56 72 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 72 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 72 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 60 72 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 59 72 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 59 72 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 72 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 72 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 58 72 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 57 72 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 57 72 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 72 56 72 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 60 71 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 60 71 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 60 71 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 59 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 59 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 58 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 58 71 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 58 71 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 57 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 57 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 56 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 60 71 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 60 71 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 60 71 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 59 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 59 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 58 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 58 71 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 58 71 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 57 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 57 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 71 56 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 71 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 71 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 71 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 59 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 59 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 71 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 71 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 71 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 57 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 57 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 56 71 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 70 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 70 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 70 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 59 70 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 59 70 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 70 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 70 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 70 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 57 70 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 57 70 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 56 70 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 70 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 70 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 60 70 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 59 70 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 59 70 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 70 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 70 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 58 70 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 57 70 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 57 70 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 70 56 70 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 60 69 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 60 69 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 60 69 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 59 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 59 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 58 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 58 69 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 58 69 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 57 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 57 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 56 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 60 69 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 60 69 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 60 69 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 59 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 59 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 58 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 58 69 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 58 69 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 57 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 57 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 69 56 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 69 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 69 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 69 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 59 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 59 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 69 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 69 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 69 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 57 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 57 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 56 69 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 68 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 68 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 68 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 59 68 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 59 68 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 68 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 68 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 68 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 57 68 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 57 68 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 56 68 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 68 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 68 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 60 68 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 59 68 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 59 68 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 68 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 68 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 58 68 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 57 68 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 57 68 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 68 56 68 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 60 67 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 60 67 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 60 67 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 59 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 59 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 58 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 58 67 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 58 67 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 57 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 57 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 56 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 60 67 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 60 67 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 60 67 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 59 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 59 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 58 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 58 67 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 58 67 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 57 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 57 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 67 56 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 60 67 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 60 67 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 60 67 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 59 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 59 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 58 67 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 58 67 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 58 67 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 57 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 57 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 56 67 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 60 66 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 60 66 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 60 66 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 59 66 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 59 66 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 58 66 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 58 66 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 58 66 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 57 66 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 57 66 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 66 56 66 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 66 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 66 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 66 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 59 66 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 59 66 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 66 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 66 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 66 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 57 66 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 57 66 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 56 66 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 65 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 65 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 65 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 59 65 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 59 65 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 65 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 65 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 65 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 57 65 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 57 65 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 56 65 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 65 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 65 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 60 65 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 59 65 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 59 65 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 65 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 65 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 58 65 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 57 65 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 57 65 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 65 56 65 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 60 64 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 60 64 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 60 64 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 59 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 59 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 58 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 58 64 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 58 64 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 57 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 57 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 56 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 60 64 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 60 64 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 60 64 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 59 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 59 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 58 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 58 64 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 58 64 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 57 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 57 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 64 56 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 64 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 64 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 64 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 59 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 59 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 64 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 64 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 64 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 57 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 57 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 56 64 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 63 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 63 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 63 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 59 63 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 59 63 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 63 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 63 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 63 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 57 63 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 57 63 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 56 63 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 63 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 63 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 60 63 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 59 63 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 59 63 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 63 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 63 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 58 63 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 57 63 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 57 63 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 63 56 63 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 60 62 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 60 62 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 60 62 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 59 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 59 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 58 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 58 62 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 58 62 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 57 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 57 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 56 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 60 62 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 60 62 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 60 62 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 59 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 59 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 58 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 58 62 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 58 62 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 57 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 57 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 62 56 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 62 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 62 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 62 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 59 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 59 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 62 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 62 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 62 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 57 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 57 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 56 62 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 61 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 61 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 61 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 59 61 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 59 61 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 61 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 61 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 61 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 57 61 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 57 61 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 56 61 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 61 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 61 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 60 61 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 59 61 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 59 61 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 61 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 61 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 58 61 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 57 61 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 57 61 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 61 56 61 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 60 60 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 60 60 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 60 60 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 59 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 59 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 58 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 58 60 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 58 60 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 57 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 57 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 56 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 60 60 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 60 60 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 60 60 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 59 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 59 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 58 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 58 60 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 58 60 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 57 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 57 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 60 56 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 60 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 60 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 60 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 59 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 59 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 60 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 60 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 60 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 57 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 57 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 56 60 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 59 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 59 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 59 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 59 59 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 59 59 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 59 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 59 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 59 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 57 59 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 57 59 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 56 59 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 59 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 59 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 60 59 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 59 59 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 59 59 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 59 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 59 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 58 59 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 57 59 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 57 59 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 59 56 59 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 60 58 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 60 58 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 60 58 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 59 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 59 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 58 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 58 58 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 58 58 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 57 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 57 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 56 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 60 58 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 60 58 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 60 58 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 59 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 59 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 58 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 58 58 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 58 58 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 57 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 57 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 58 56 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 58 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 58 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 58 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 59 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 59 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 58 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 58 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 58 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 57 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 57 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 56 58 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 57 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 57 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 57 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 59 57 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 59 57 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 57 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 57 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 57 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 57 57 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 57 57 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 56 57 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 57 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 57 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 60 57 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 59 57 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 59 57 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 57 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 57 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 58 57 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 57 57 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 57 57 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 57 56 57 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 60 56 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 60 56 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 60 56 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 59 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 59 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 58 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 58 56 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 58 56 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 57 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 57 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 56 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 60 56 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 60 56 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 60 56 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 59 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 59 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 58 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 58 56 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 58 56 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 57 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 57 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 56 56 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 56 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 56 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 56 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 59 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 59 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 56 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 56 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 56 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 57 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 57 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 56 56 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 55 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 55 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 55 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 59 55 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 59 55 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 55 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 55 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 55 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 57 55 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 57 55 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 56 55 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 55 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 55 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 60 55 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 59 55 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 59 55 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 55 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 55 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 58 55 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 57 55 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 57 55 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 55 56 55 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 60 54 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 60 54 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 60 54 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 59 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 59 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 58 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 58 54 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 58 54 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 57 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 57 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 56 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 60 54 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 60 54 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 60 54 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 59 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 59 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 58 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 58 54 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 58 54 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 57 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 57 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 54 56 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 60 54 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 60 54 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 60 54 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 59 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 59 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 58 54 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 58 54 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 58 54 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 57 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 57 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 56 54 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 60 53 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 60 53 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 60 53 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 59 53 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 59 53 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 58 53 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 58 53 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 58 53 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 57 53 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 57 53 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 53 56 53 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 53 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 53 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 53 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 59 53 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 59 53 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 53 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 53 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 53 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 57 53 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 57 53 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 56 53 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 52 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 52 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 52 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 59 52 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 59 52 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 52 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 52 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 52 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 57 52 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 57 52 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 56 52 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 52 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 52 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 60 52 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 59 52 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 59 52 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 52 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 52 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 58 52 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 57 52 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 57 52 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 52 56 52 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 60 51 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 60 51 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 60 51 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 59 51 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 59 51 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 58 51 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 58 51 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 58 51 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 57 51 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 57 51 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 56 51 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 60 51 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 60 51 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 60 51 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 59 51 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 59 51 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 58 51 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 58 51 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 58 51 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 57 51 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 57 51 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 51 56 51 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 60 24 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 60 24 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 60 24 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 59 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 59 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 58 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 58 24 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 58 24 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 57 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 57 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 56 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 60 24 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 60 24 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 60 24 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 59 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 59 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 58 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 58 24 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 58 24 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 57 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 57 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 24 56 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 60 24 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 60 24 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 60 24 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 59 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 59 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 58 24 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 58 24 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 58 24 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 57 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 57 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 56 24 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 60 23 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 60 23 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 60 23 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 59 23 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 59 23 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 58 23 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 58 23 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 58 23 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 57 23 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 57 23 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 23 56 23 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 23 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 23 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 23 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 59 23 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 59 23 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 23 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 23 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 23 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 57 23 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 57 23 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 56 23 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 22 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 22 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 22 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 59 22 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 59 22 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 22 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 22 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 22 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 57 22 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 57 22 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 56 22 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 22 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 22 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 60 22 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 59 22 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 59 22 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 22 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 22 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 58 22 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 57 22 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 57 22 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 22 56 22 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 60 21 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 60 21 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 60 21 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 59 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 59 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 58 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 58 21 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 58 21 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 57 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 57 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 56 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 60 21 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 60 21 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 60 21 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 59 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 59 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 58 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 58 21 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 58 21 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 57 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 57 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 21 56 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 21 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 21 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 21 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 59 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 59 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 21 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 21 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 21 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 57 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 57 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 56 21 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 20 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 20 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 20 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 59 20 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 59 20 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 20 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 20 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 20 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 57 20 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 57 20 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 56 20 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 20 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 20 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 60 20 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 59 20 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 59 20 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 20 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 20 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 58 20 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 57 20 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 57 20 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 20 56 20 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 60 19 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 60 19 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 60 19 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 59 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 59 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 58 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 58 19 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 58 19 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 57 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 57 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 56 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 60 19 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 60 19 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 60 19 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 59 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 59 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 58 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 58 19 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 58 19 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 57 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 57 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 19 56 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 19 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 19 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 19 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 59 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 59 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 19 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 19 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 19 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 57 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 57 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 56 19 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 18 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 18 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 18 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 59 18 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 59 18 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 18 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 18 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 18 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 57 18 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 57 18 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 56 18 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 18 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 18 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 60 18 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 59 18 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 59 18 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 18 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 18 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 58 18 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 57 18 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 57 18 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 18 56 18 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 60 17 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 60 17 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 60 17 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 59 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 59 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 58 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 58 17 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 58 17 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 57 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 57 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 56 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 60 17 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 60 17 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 60 17 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 59 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 59 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 58 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 58 17 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 58 17 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 57 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 57 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 17 56 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 17 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 17 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 17 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 59 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 59 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 17 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 17 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 17 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 57 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 57 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 56 17 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 16 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 16 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 16 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 59 16 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 59 16 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 16 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 16 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 16 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 57 16 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 57 16 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 56 16 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 16 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 16 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 60 16 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 59 16 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 59 16 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 16 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 16 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 58 16 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 57 16 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 57 16 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 16 56 16 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 60 15 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 60 15 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 60 15 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 59 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 59 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 58 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 58 15 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 58 15 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 57 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 57 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 56 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 60 15 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 60 15 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 60 15 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 59 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 59 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 58 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 58 15 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 58 15 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 57 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 57 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 15 56 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 15 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 15 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 15 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 59 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 59 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 15 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 15 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 15 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 57 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 57 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 56 15 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 14 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 14 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 14 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 59 14 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 59 14 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 14 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 14 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 14 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 57 14 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 57 14 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 56 14 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 14 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 14 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 60 14 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 59 14 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 59 14 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 14 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 14 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 58 14 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 57 14 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 57 14 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 14 56 14 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 60 13 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 60 13 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 60 13 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 59 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 59 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 58 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 58 13 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 58 13 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 57 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 57 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 56 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 60 13 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 60 13 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 60 13 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 59 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 59 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 58 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 58 13 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 58 13 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 57 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 57 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 13 56 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 13 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 13 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 13 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 59 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 59 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 13 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 13 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 13 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 57 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 57 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 56 13 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 12 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 12 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 12 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 59 12 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 59 12 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 12 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 12 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 12 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 57 12 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 57 12 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 56 12 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 12 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 12 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 60 12 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 59 12 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 59 12 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 12 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 12 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 58 12 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 57 12 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 57 12 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 12 56 12 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 60 11 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 60 11 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 60 11 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 59 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 59 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 58 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 58 11 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 58 11 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 57 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 57 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 56 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 60 11 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 60 11 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 60 11 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 59 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 59 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 58 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 58 11 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 58 11 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 57 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 57 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 11 56 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 11 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 11 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 11 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 59 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 59 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 11 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 11 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 11 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 57 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 57 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 56 11 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 10 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 10 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 10 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 59 10 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 59 10 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 10 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 10 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 10 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 57 10 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 57 10 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 56 10 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 10 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 10 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 60 10 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 59 10 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 59 10 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 10 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 10 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 58 10 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 57 10 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 57 10 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 10 56 10 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 60 9 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 60 9 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 60 9 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 59 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 59 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 58 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 58 9 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 58 9 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 57 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 57 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 56 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 60 9 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 60 9 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 60 9 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 59 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 59 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 58 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 58 9 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 58 9 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 57 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 57 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 9 56 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 9 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 9 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 9 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 59 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 59 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 9 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 9 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 9 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 57 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 57 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 56 9 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 8 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 8 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 8 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 59 8 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 59 8 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 8 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 8 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 8 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 57 8 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 57 8 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 56 8 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 8 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 8 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 60 8 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 59 8 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 59 8 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 8 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 8 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 58 8 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 57 8 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 57 8 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 8 56 8 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 60 7 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 60 7 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 60 7 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 59 7 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 59 7 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 58 7 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 58 7 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 58 7 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 57 7 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 57 7 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 56 7 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 60 7 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 60 7 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 60 7 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 59 7 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 59 7 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 58 7 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 58 7 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 58 7 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 57 7 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 57 7 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 7 56 7 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 60 6 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 60 6 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 60 6 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 59 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 59 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 58 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 58 6 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 58 6 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 57 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 57 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 56 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 60 6 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 60 6 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 60 6 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 59 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 59 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 58 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 58 6 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 58 6 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 57 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 57 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 6 56 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 6 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 6 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 6 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 59 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 59 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 6 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 6 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 6 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 57 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 57 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 56 6 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 5 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 5 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 5 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 59 5 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 59 5 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 5 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 5 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 5 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 57 5 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 57 5 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 56 5 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 5 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 5 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 60 5 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 59 5 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 59 5 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 5 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 5 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 58 5 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 57 5 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 57 5 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 5 56 5 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 60 4 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 60 4 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 60 4 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 59 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 59 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 58 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 58 4 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 58 4 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 57 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 57 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 56 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 60 4 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 60 4 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 60 4 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 59 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 59 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 58 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 58 4 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 58 4 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 57 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 57 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 4 56 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 4 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 4 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 4 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 59 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 59 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 4 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 4 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 4 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 57 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 57 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 56 4 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 3 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 3 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 3 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 59 3 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 59 3 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 3 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 3 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 3 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 57 3 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 57 3 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 56 3 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 3 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 3 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 60 3 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 59 3 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 59 3 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 3 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 3 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 58 3 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 57 3 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 57 3 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 3 56 3 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 60 2 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 60 2 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 60 2 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 59 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 59 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 58 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 58 2 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 58 2 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 57 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 57 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 56 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 60 2 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 60 2 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 60 2 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 59 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 59 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 58 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 58 2 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 58 2 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 57 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 57 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 2 56 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 2 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 2 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 2 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 59 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 59 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 2 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 2 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 2 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 57 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 57 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 56 2 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 1 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 1 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 1 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 59 1 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 59 1 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 1 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 1 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 1 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 57 1 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 57 1 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 56 1 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 1 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 1 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 60 1 60 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 59 1 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 59 1 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 1 59 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 1 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 58 1 58 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 57 1 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 57 1 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel nfet_brown s 1 56 1 57 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 198
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
