magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 8 0 8 7 6 C0
port 1 nsew
rlabel  s 7 0 7 7 6 C0
port 1 nsew
rlabel  s 6 0 7 7 6 C0
port 1 nsew
rlabel  s 6 0 6 7 6 C0
port 1 nsew
rlabel  s 5 0 5 7 6 C0
port 1 nsew
rlabel  s 5 0 5 7 6 C0
port 1 nsew
rlabel  s 4 0 4 7 6 C0
port 1 nsew
rlabel  s 4 0 4 7 6 C0
port 1 nsew
rlabel  s 3 0 3 7 6 C0
port 1 nsew
rlabel  s 3 0 3 7 6 C0
port 1 nsew
rlabel  s 2 0 2 7 6 C0
port 1 nsew
rlabel  s 1 0 2 7 6 C0
port 1 nsew
rlabel  s 1 0 1 7 6 C0
port 1 nsew
rlabel  s 0 0 0 7 4 C0
port 1 nsew
rlabel  s 0 0 0 7 4 C0
port 1 nsew
rlabel  s 0 0 8 0 8 C0
port 1 nsew
rlabel  s 8 0 8 8 6 C1
port 2 nsew
rlabel  s 7 0 7 8 6 C1
port 2 nsew
rlabel  s 7 0 7 8 6 C1
port 2 nsew
rlabel  s 6 0 6 8 6 C1
port 2 nsew
rlabel  s 6 0 6 8 6 C1
port 2 nsew
rlabel  s 5 0 5 8 6 C1
port 2 nsew
rlabel  s 4 0 5 8 6 C1
port 2 nsew
rlabel  s 4 0 4 8 6 C1
port 2 nsew
rlabel  s 3 0 4 8 6 C1
port 2 nsew
rlabel  s 3 0 3 8 6 C1
port 2 nsew
rlabel  s 2 0 2 8 6 C1
port 2 nsew
rlabel  s 2 0 2 8 6 C1
port 2 nsew
rlabel  s 1 0 1 8 6 C1
port 2 nsew
rlabel  s 1 0 1 8 6 C1
port 2 nsew
rlabel  s 0 0 0 8 4 C1
port 2 nsew
rlabel  s 0 8 8 8 6 C1
port 2 nsew
rlabel metal_blue s 4 4 4 4 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 9 8
string LEFview TRUE
<< end >>
