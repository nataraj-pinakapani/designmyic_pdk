magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel � s 50 -2 74 24 6 DRN_HVC
port 3 nsew power bidirectional
rlabel 
 s 38 -2 49 10 6 DRN_HVC
port 3 nsew power bidirectional
rlabel � s 0 -2 24 0 8 SRC_BDY_HVC
port 4 nsew ground bidirectional
rlabel 
 s 26 -2 37 10 6 SRC_BDY_HVC
port 4 nsew ground bidirectional
rlabel  s 7 103 68 164 6 VSSIO_PAD
port 5 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 6 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 6 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 54 75 55 6 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 46 75 46 6 VSSA
port 6 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 6 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 6 nsew ground bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 7 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 7 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 7 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 7 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 8 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 8 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 8 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 8 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 9 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 9 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 9 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 9 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 10 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 10 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 10 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 10 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 12 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 12 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 12 nsew power bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 12 nsew power bidirectional
rlabel  s 1 190 1 190 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 13 nsew ground bidirectional
rlabel 
 s 0 -2 24 24 6 VSSIO
port 13 nsew ground bidirectional
rlabel 
 s 50 -2 74 24 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 13 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 14 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 14 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 14 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 14 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 15 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 15 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 15 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 15 nsew ground bidirectional
<< properties >>
string LEFclass PAD POWER
string FIXED_BBOX 0 0 75 198
string LEFview TRUE
<< end >>
