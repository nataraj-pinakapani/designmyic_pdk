magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 3 10 5 6 DRAIN
port 1 nsew
rlabel  s 1 6 9 6 6 GATE
port 2 nsew
rlabel  s 1 0 9 0 8 GATE
port 2 nsew
rlabel  s 0 1 10 3 6 SOURCE
port 3 nsew
rlabel  s 0 1 0 5 4 SUBSTRATE
port 4 nsew
rlabel  s 9 1 10 5 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 10 6
string LEFview TRUE
<< end >>
