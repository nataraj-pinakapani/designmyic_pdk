magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal default
rlabel  s 74 53 75 56 6 AMUXBUS_A
port 1 nsew signal default
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal default
rlabel  s 74 48 75 51 6 AMUXBUS_B
port 2 nsew signal default
rlabel  s 0 9 1 14 4 VCCD
port 3 nsew signal default
rlabel  s 74 9 75 14 6 VCCD
port 3 nsew signal default
rlabel  s 0 9 1 13 4 VCCD
port 3 nsew signal default
rlabel  s 74 9 75 13 6 VCCD
port 3 nsew signal default
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew signal default
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew signal default
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew signal default
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew signal default
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew signal default
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew signal default
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew signal default
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew signal default
rlabel  s 0 20 24 24 6 VDDIO
port 6 nsew signal default
rlabel  s 0 95 1 95 4 VDDIO
port 6 nsew signal default
rlabel  s 0 91 20 95 6 VDDIO
port 6 nsew signal default
rlabel  s 0 90 1 91 4 VDDIO
port 6 nsew signal default
rlabel  s 0 70 24 90 6 VDDIO
port 6 nsew signal default
rlabel  s 0 70 1 70 4 VDDIO
port 6 nsew signal default
rlabel  s 50 20 75 24 6 VDDIO
port 6 nsew signal default
rlabel  s 74 95 75 95 6 VDDIO
port 6 nsew signal default
rlabel  s 74 90 75 91 6 VDDIO
port 6 nsew signal default
rlabel  s 74 70 75 70 6 VDDIO
port 6 nsew signal default
rlabel  s 55 91 75 95 6 VDDIO
port 6 nsew signal default
rlabel  s 51 70 75 90 6 VDDIO
port 6 nsew signal default
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew signal default
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew signal default
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew signal default
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew signal default
rlabel  s 0 64 24 69 6 VDDIO_Q
port 7 nsew signal default
rlabel  s 50 64 75 69 6 VDDIO_Q
port 7 nsew signal default
rlabel  s 0 64 1 68 4 VDDIO_Q
port 7 nsew signal default
rlabel  s 74 64 75 68 6 VDDIO_Q
port 7 nsew signal default
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew signal default
rlabel  s 0 48 1 48 4 VSSA
port 8 nsew signal default
rlabel  s 0 52 1 53 4 VSSA
port 8 nsew signal default
rlabel  s 0 56 1 57 4 VSSA
port 8 nsew signal default
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew signal default
rlabel  s 74 48 75 48 6 VSSA
port 8 nsew signal default
rlabel  s 74 52 75 53 6 VSSA
port 8 nsew signal default
rlabel  s 74 56 75 57 6 VSSA
port 8 nsew signal default
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew signal default
rlabel  s 0 48 1 57 4 VSSA
port 8 nsew signal default
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew signal default
rlabel  s 74 48 75 57 6 VSSA
port 8 nsew signal default
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew signal default
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew signal default
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew signal default
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew signal default
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew signal default
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew signal default
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew signal default
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew signal default
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew signal default
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew signal default
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew signal default
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew signal default
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew signal default
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew signal default
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew signal default
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew signal default
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew signal default
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew signal default
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew signal default
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew signal default
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
