/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/xschem/xschem_verilog_import/spm.spice