magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 139 53 140 56 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 139 48 140 51 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel 
 s 8 14 9 14 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 8 14 8 14 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 8 14 8 14 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 8 0 8 14 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 8 14 9 14 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 8 14 9 14 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 8 14 9 14 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 65 1 66 1 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 65 0 66 1 8 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 65 1 66 1 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 65 1 66 1 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 52 8 52 8 6 ANALOG_SEL
port 5 nsew signal input
rlabel 
 s 52 8 52 8 6 ANALOG_SEL
port 5 nsew signal input
rlabel 
 s 52 8 52 8 6 ANALOG_SEL
port 5 nsew signal input
rlabel 
 s 52 0 52 8 6 ANALOG_SEL
port 5 nsew signal input
rlabel 
 s 129 0 129 21 6 DM[0]
port 6 nsew signal input
rlabel 
 s 129 21 129 22 6 DM[0]
port 6 nsew signal input
rlabel 
 s 128 20 129 22 6 DM[1]
port 7 nsew signal input
rlabel 
 s 128 20 129 20 6 DM[1]
port 7 nsew signal input
rlabel 
 s 128 20 129 20 6 DM[1]
port 7 nsew signal input
rlabel 
 s 128 20 129 20 6 DM[1]
port 7 nsew signal input
rlabel 
 s 128 20 129 20 6 DM[1]
port 7 nsew signal input
rlabel 
 s 128 20 129 20 6 DM[1]
port 7 nsew signal input
rlabel 
 s 128 0 129 20 6 DM[1]
port 7 nsew signal input
rlabel 
 s 108 0 109 20 6 DM[2]
port 8 nsew signal input
rlabel 
 s 108 21 109 22 6 DM[2]
port 8 nsew signal input
rlabel 
 s 108 20 109 21 6 DM[2]
port 8 nsew signal input
rlabel 
 s 22 32 23 32 6 ENABLE_H
port 9 nsew signal input
rlabel 
 s 22 32 23 32 6 ENABLE_H
port 9 nsew signal input
rlabel 
 s 22 32 22 32 6 ENABLE_H
port 9 nsew signal input
rlabel 
 s 22 0 22 32 6 ENABLE_H
port 9 nsew signal input
rlabel 
 s 7 0 7 20 6 ENABLE_INP_H
port 10 nsew signal input
rlabel 
 s 9 0 9 9 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel 
 s 96 0 96 2 6 ENABLE_VDDIO
port 12 nsew signal input
rlabel 
 s 6 0 6 13 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel 
 s 20 18 20 23 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 18 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 20 0 20 18 6 HLD_H_N
port 14 nsew signal input
rlabel 
 s 27 14 28 14 6 HLD_OVR
port 15 nsew signal input
rlabel 
 s 27 0 28 14 6 HLD_OVR
port 15 nsew signal input
rlabel 
 s 27 14 28 14 6 HLD_OVR
port 15 nsew signal input
rlabel 
 s 27 14 28 14 6 HLD_OVR
port 15 nsew signal input
rlabel 
 s 27 14 28 14 6 HLD_OVR
port 15 nsew signal input
rlabel 
 s 27 14 28 14 6 HLD_OVR
port 15 nsew signal input
rlabel 
 s 45 8 46 8 6 HYS_TRIM
port 16 nsew signal input
rlabel 
 s 45 0 46 8 6 HYS_TRIM
port 16 nsew signal input
rlabel 
 s 45 8 46 8 6 HYS_TRIM
port 16 nsew signal input
rlabel 
 s 45 8 46 8 6 HYS_TRIM
port 16 nsew signal input
rlabel 
 s 45 8 46 8 6 HYS_TRIM
port 16 nsew signal input
rlabel 
 s 87 0 87 22 6 IB_MODE_SEL[0]
port 17 nsew signal input
rlabel 
 s 67 0 67 22 6 IB_MODE_SEL[1]
port 18 nsew signal input
rlabel 
 s 20 0 21 15 6 IN
port 19 nsew signal output
rlabel 
 s 108 8 108 8 6 INP_DIS
port 20 nsew signal input
rlabel 
 s 108 0 108 8 6 INP_DIS
port 20 nsew signal input
rlabel 
 s 107 8 108 8 6 INP_DIS
port 20 nsew signal input
rlabel 
 s 107 8 108 8 6 INP_DIS
port 20 nsew signal input
rlabel 
 s 107 8 108 8 6 INP_DIS
port 20 nsew signal input
rlabel 
 s 24 0 25 0 8 IN_H
port 21 nsew signal output
rlabel 
 s 24 0 25 0 8 IN_H
port 21 nsew signal output
rlabel 
 s 24 0 25 1 8 IN_H
port 21 nsew signal output
rlabel 
 s 24 1 25 1 6 IN_H
port 21 nsew signal output
rlabel 
 s 23 1 25 1 6 IN_H
port 21 nsew signal output
rlabel 
 s 124 8 125 8 6 OE_N
port 22 nsew signal input
rlabel 
 s 124 0 125 8 6 OE_N
port 22 nsew signal input
rlabel 
 s 124 8 125 8 6 OE_N
port 22 nsew signal input
rlabel 
 s 124 8 125 8 6 OE_N
port 22 nsew signal input
rlabel 
 s 78 34 79 51 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 79 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 31 79 31 6 OUT
port 23 nsew signal input
rlabel 
 s 78 15 79 31 6 OUT
port 23 nsew signal input
rlabel 
 s 78 15 79 15 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 79 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 31 79 31 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 79 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 15 79 15 6 OUT
port 23 nsew signal input
rlabel 
 s 78 31 79 31 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 78 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 31 78 31 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 78 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 31 78 31 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 78 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 78 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 34 78 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 32 78 34 6 OUT
port 23 nsew signal input
rlabel 
 s 78 32 78 32 6 OUT
port 23 nsew signal input
rlabel 
 s 78 32 78 32 6 OUT
port 23 nsew signal input
rlabel 
 s 78 31 78 32 6 OUT
port 23 nsew signal input
rlabel 
 s 78 15 79 15 6 OUT
port 23 nsew signal input
rlabel 
 s 78 51 79 51 6 OUT
port 23 nsew signal input
rlabel 
 s 74 15 79 15 6 OUT
port 23 nsew signal input
rlabel 
 s 74 14 75 15 6 OUT
port 23 nsew signal input
rlabel 
 s 74 14 75 14 6 OUT
port 23 nsew signal input
rlabel 
 s 74 14 74 14 6 OUT
port 23 nsew signal input
rlabel 
 s 74 0 74 14 6 OUT
port 23 nsew signal input
rlabel  s 40 133 63 148 6 PAD
port 24 nsew signal bidirectional
rlabel 
 s 4 74 5 160 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 4 74 5 74 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 4 73 5 74 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 4 73 5 73 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 4 73 5 73 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 4 73 4 73 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 73 4 73 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 73 4 73 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 73 4 73 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 72 4 73 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 72 4 72 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 72 3 72 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 72 3 72 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 72 3 72 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 72 3 72 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 72 3 72 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 71 3 72 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 71 3 71 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 71 2 71 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 5 2 5 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 0 2 5 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 2 71 2 71 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 5 2 5 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 71 2 71 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 5 2 5 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 71 2 71 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 71 2 71 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 6 2 71 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 6 2 6 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 6 2 6 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 5 2 6 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 1 5 2 5 6 PAD_A_ESD_0_H
port 25 nsew signal bidirectional
rlabel 
 s 3 74 4 161 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 3 74 4 74 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 3 74 4 74 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 3 74 3 74 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 3 73 3 74 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 2 73 3 73 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 2 73 3 73 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 2 73 3 73 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 2 73 3 73 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 2 73 3 73 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 2 73 2 73 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 2 72 2 73 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 1 72 2 72 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 1 72 2 72 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 1 72 2 72 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 1 72 2 72 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 1 72 2 72 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 1 72 1 72 6 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 0 71 1 72 4 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 0 71 1 71 4 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 0 71 1 71 4 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 0 0 1 71 4 PAD_A_ESD_1_H
port 26 nsew signal bidirectional
rlabel 
 s 5 73 6 123 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 5 73 6 73 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 5 73 6 73 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 5 73 5 73 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 5 73 5 73 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 4 72 5 73 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 4 72 5 72 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 4 72 5 72 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 4 72 5 72 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 4 72 5 72 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 4 72 4 72 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 4 72 4 72 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 71 4 72 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 71 4 71 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 71 4 71 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 71 4 71 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 6 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 0 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 71 3 71 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 6 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 71 3 71 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 6 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 3 6 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 71 3 71 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 6 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 70 3 71 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 6 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 70 3 70 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 70 3 70 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 7 3 70 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 7 3 7 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 6 3 7 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 2 6 3 6 6 PAD_A_NOESD_H
port 27 nsew signal bidirectional
rlabel 
 s 66 0 66 22 6 SLEW_CTL[0]
port 28 nsew signal input
rlabel 
 s 46 0 47 22 6 SLEW_CTL[1]
port 29 nsew signal input
rlabel 
 s 125 19 125 31 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 0 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 19 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 18 125 19 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 13 125 18 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 13 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 125 12 125 12 6 SLOW
port 30 nsew signal input
rlabel 
 s 131 110 131 110 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 131 62 131 110 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 131 62 131 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 131 110 131 110 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 131 62 131 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 131 62 131 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 131 62 131 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 130 110 131 111 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 130 62 131 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 130 62 131 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 130 62 130 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 130 62 130 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 130 61 130 62 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 130 0 130 61 6 TIE_HI_ESD
port 31 nsew signal output
rlabel 
 s 115 111 116 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 0 116 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 111 116 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 111 116 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 111 116 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 111 116 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 111 116 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 111 115 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 115 111 115 111 6 TIE_LO_ESD
port 32 nsew signal output
rlabel 
 s 44 5 45 5 6 VINREF
port 33 nsew signal input
rlabel 
 s 44 5 45 5 6 VINREF
port 33 nsew signal input
rlabel 
 s 44 5 45 5 6 VINREF
port 33 nsew signal input
rlabel 
 s 44 4 44 5 6 VINREF
port 33 nsew signal input
rlabel 
 s 44 0 44 4 6 VINREF
port 33 nsew signal input
rlabel 
 s 88 0 88 22 6 VTRIP_SEL
port 34 nsew signal input
rlabel  s 0 9 1 14 4 VCCD
port 35 nsew power bidirectional
rlabel  s 139 13 140 14 6 VCCD
port 35 nsew power bidirectional
rlabel  s 139 9 140 9 6 VCCD
port 35 nsew power bidirectional
rlabel  s 138 9 140 13 6 VCCD
port 35 nsew power bidirectional
rlabel  s 0 9 1 13 4 VCCD
port 35 nsew power bidirectional
rlabel  s 139 9 140 13 6 VCCD
port 35 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 36 nsew power bidirectional
rlabel  s 139 2 140 7 6 VCCHIB
port 36 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 36 nsew power bidirectional
rlabel  s 139 2 140 7 6 VCCHIB
port 36 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 37 nsew power bidirectional
rlabel  s 139 15 140 18 6 VDDA
port 37 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 37 nsew power bidirectional
rlabel  s 139 15 140 18 6 VDDA
port 37 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 38 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 38 nsew power bidirectional
rlabel  s 139 20 140 24 6 VDDIO
port 38 nsew power bidirectional
rlabel  s 139 70 140 95 6 VDDIO
port 38 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 38 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 38 nsew power bidirectional
rlabel  s 139 20 140 24 6 VDDIO
port 38 nsew power bidirectional
rlabel  s 139 70 140 95 6 VDDIO
port 38 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 39 nsew power bidirectional
rlabel  s 139 64 140 69 6 VDDIO_Q
port 39 nsew power bidirectional
rlabel  s 0 64 1 68 4 VDDIO_Q
port 39 nsew power bidirectional
rlabel  s 139 64 140 68 6 VDDIO_Q
port 39 nsew power bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 40 nsew ground bidirectional
rlabel  s 0 48 1 48 4 VSSA
port 40 nsew ground bidirectional
rlabel  s 0 52 1 53 4 VSSA
port 40 nsew ground bidirectional
rlabel  s 0 56 1 57 4 VSSA
port 40 nsew ground bidirectional
rlabel  s 139 37 140 40 6 VSSA
port 40 nsew ground bidirectional
rlabel  s 139 48 140 48 6 VSSA
port 40 nsew ground bidirectional
rlabel  s 139 52 140 53 6 VSSA
port 40 nsew ground bidirectional
rlabel  s 139 56 140 57 6 VSSA
port 40 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 40 nsew ground bidirectional
rlabel  s 0 48 1 57 4 VSSA
port 40 nsew ground bidirectional
rlabel  s 139 37 140 40 6 VSSA
port 40 nsew ground bidirectional
rlabel  s 139 48 140 57 6 VSSA
port 40 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 41 nsew ground bidirectional
rlabel  s 139 42 140 46 6 VSSD
port 41 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 41 nsew ground bidirectional
rlabel  s 139 42 140 46 6 VSSD
port 41 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 42 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 42 nsew ground bidirectional
rlabel  s 139 176 140 200 6 VSSIO
port 42 nsew ground bidirectional
rlabel  s 139 26 140 30 6 VSSIO
port 42 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 42 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 42 nsew ground bidirectional
rlabel  s 139 176 140 200 6 VSSIO
port 42 nsew ground bidirectional
rlabel  s 139 26 140 30 6 VSSIO
port 42 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 43 nsew ground bidirectional
rlabel  s 139 58 140 63 6 VSSIO_Q
port 43 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 43 nsew ground bidirectional
rlabel  s 139 58 140 63 6 VSSIO_Q
port 43 nsew ground bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 44 nsew power bidirectional
rlabel  s 139 32 140 35 6 VSWITCH
port 44 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 44 nsew power bidirectional
rlabel  s 139 32 140 35 6 VSWITCH
port 44 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 140 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
