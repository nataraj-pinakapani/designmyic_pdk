magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 1 1 2 2 6 DRAIN
port 1 nsew
rlabel  s 1 2 2 2 6 DRAIN
port 1 nsew
rlabel  s 1 1 1 2 6 DRAIN
port 1 nsew
rlabel  s 0 2 2 3 6 GATE
port 2 nsew
rlabel  s 2 0 2 2 6 SOURCE
port 3 nsew
rlabel  s 1 0 1 2 6 SOURCE
port 3 nsew
rlabel  s 0 0 0 2 4 SOURCE
port 3 nsew
rlabel  s 0 0 2 0 8 SOURCE
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 2 3
string LEFview TRUE
<< end >>
