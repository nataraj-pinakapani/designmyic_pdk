magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 2 4 4 6 DRAIN
port 1 nsew
rlabel  s 1 6 4 6 6 GATE
port 2 nsew
rlabel  s 1 0 4 0 8 GATE
port 2 nsew
rlabel  s 0 4 4 6 6 SOURCE
port 3 nsew
rlabel  s 0 1 4 2 6 SOURCE
port 3 nsew
rlabel  s 0 1 0 6 4 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 4 6
string LEFview TRUE
<< end >>
