magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 6 0 7 6 6 C0
port 1 nsew
rlabel  s 5 4 6 6 6 C0
port 1 nsew
rlabel  s 5 0 6 3 6 C0
port 1 nsew
rlabel  s 4 4 4 6 6 C0
port 1 nsew
rlabel  s 4 0 4 3 6 C0
port 1 nsew
rlabel  s 3 4 3 6 6 C0
port 1 nsew
rlabel  s 3 0 3 3 6 C0
port 1 nsew
rlabel  s 1 4 2 6 6 C0
port 1 nsew
rlabel  s 1 0 2 3 6 C0
port 1 nsew
rlabel  s 0 6 7 6 6 C0
port 1 nsew
rlabel  s 0 0 0 6 4 C0
port 1 nsew
rlabel  s 0 0 7 0 8 C0
port 1 nsew
rlabel  s 6 3 6 5 6 C1
port 2 nsew
rlabel  s 6 1 6 3 6 C1
port 2 nsew
rlabel  s 5 3 5 5 6 C1
port 2 nsew
rlabel  s 5 1 5 3 6 C1
port 2 nsew
rlabel  s 3 3 4 5 6 C1
port 2 nsew
rlabel  s 3 1 4 3 6 C1
port 2 nsew
rlabel  s 2 3 2 5 6 C1
port 2 nsew
rlabel  s 2 1 2 3 6 C1
port 2 nsew
rlabel  s 1 3 1 5 6 C1
port 2 nsew
rlabel  s 1 3 6 3 6 C1
port 2 nsew
rlabel  s 1 1 1 3 6 C1
port 2 nsew
rlabel  s 0 0 7 6 6 MET4
port 3 nsew
rlabel metal_blue s 3 4 3 5 6 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 7 6
string LEFview TRUE
<< end >>
