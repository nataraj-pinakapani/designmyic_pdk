magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< dnwell >>
rect 0 4453 7789 4845
rect 0 3943 12122 4453
rect 0 1679 12172 3943
rect 0 766 12061 1679
rect 7592 659 12061 766
rect 10479 545 12061 659
<< nwell >>
rect 9756 4966 10366 4968
rect 7709 4925 12206 4966
rect -84 4576 12206 4925
rect -84 3937 12338 4576
rect -84 3907 10300 3937
rect -84 3560 290 3907
rect 897 3621 10300 3907
rect 1948 3589 10300 3621
rect -84 2240 206 3560
rect 1948 3476 3112 3589
rect 11966 3339 12338 3937
rect 11966 2493 12179 3339
rect -84 2024 1342 2240
rect 3110 2170 4530 2248
rect 3110 2070 5740 2170
rect 3110 2066 4530 2070
rect -84 970 702 2024
rect 9089 1604 9287 2020
rect 10088 1713 10254 2335
rect 10146 1705 10254 1713
rect 11966 1705 12493 2493
rect 11614 1090 12493 1705
rect 11614 970 12179 1090
rect -84 909 12179 970
rect -240 677 12179 909
rect -240 631 12165 677
rect -240 566 10 631
rect 10469 561 12165 631
rect 10469 541 12148 561
<< pwell >>
rect 9131 2873 9285 3525
rect 8437 1038 8723 1980
<< mvpsubdiff >>
rect 9157 3475 9259 3499
rect 9191 3441 9225 3475
rect 9157 3401 9259 3441
rect 9191 3367 9225 3401
rect 9157 3327 9259 3367
rect 9191 3293 9225 3327
rect 9157 3253 9259 3293
rect 9191 3219 9225 3253
rect 9157 3179 9259 3219
rect 9191 3145 9225 3179
rect 9157 3105 9259 3145
rect 9191 3071 9225 3105
rect 9157 3031 9259 3071
rect 9191 2997 9225 3031
rect 9157 2957 9259 2997
rect 9191 2923 9225 2957
rect 9157 2899 9259 2923
rect 8463 1930 8697 1954
rect 8497 1896 8563 1930
rect 8597 1896 8663 1930
rect 8463 1856 8697 1896
rect 8497 1822 8563 1856
rect 8597 1822 8663 1856
rect 8463 1782 8697 1822
rect 8497 1748 8563 1782
rect 8597 1748 8663 1782
rect 8463 1708 8697 1748
rect 8497 1674 8563 1708
rect 8597 1674 8663 1708
rect 8463 1634 8697 1674
rect 8497 1600 8563 1634
rect 8597 1600 8663 1634
rect 8463 1560 8697 1600
rect 8497 1526 8563 1560
rect 8597 1526 8663 1560
rect 8463 1487 8697 1526
rect 8497 1453 8563 1487
rect 8597 1453 8663 1487
rect 8463 1414 8697 1453
rect 8497 1380 8563 1414
rect 8597 1380 8663 1414
rect 8463 1341 8697 1380
rect 8497 1307 8563 1341
rect 8597 1307 8663 1341
rect 8463 1268 8697 1307
rect 8497 1234 8563 1268
rect 8597 1234 8663 1268
rect 8463 1195 8697 1234
rect 8497 1161 8563 1195
rect 8597 1161 8663 1195
rect 8463 1122 8697 1161
rect 8497 1088 8563 1122
rect 8597 1088 8663 1122
rect 8463 1064 8697 1088
<< mvnsubdiff >>
rect 7776 4858 7810 4899
rect 7844 4865 7878 4899
rect 7912 4865 7946 4899
rect 7980 4865 8014 4899
rect 8048 4865 8082 4899
rect 8116 4865 8150 4899
rect 8184 4865 8218 4899
rect 8252 4865 8286 4899
rect 8320 4865 8354 4899
rect 8388 4865 8422 4899
rect 8456 4865 8490 4899
rect 8524 4865 8558 4899
rect 8592 4865 8626 4899
rect 8660 4865 8694 4899
rect 8728 4865 8762 4899
rect 8796 4865 8830 4899
rect 8864 4865 8898 4899
rect 8932 4865 8966 4899
rect 9000 4865 9034 4899
rect 9068 4865 9102 4899
rect 9136 4865 9170 4899
rect 9204 4865 9238 4899
rect 9272 4865 9306 4899
rect 9340 4865 9374 4899
rect 9408 4865 9442 4899
rect 9476 4865 9510 4899
rect 9544 4865 9578 4899
rect 9612 4865 9646 4899
rect 9680 4865 9714 4899
rect 9748 4865 9782 4899
rect 9816 4865 9850 4899
rect 9884 4865 9918 4899
rect 9952 4865 9986 4899
rect 10020 4865 10054 4899
rect 10088 4865 10122 4899
rect 10156 4865 10190 4899
rect 10224 4865 10258 4899
rect 10292 4865 10326 4899
rect 10360 4865 10394 4899
rect 10428 4865 10462 4899
rect 10496 4865 10530 4899
rect 10564 4865 10598 4899
rect 10632 4865 10666 4899
rect 10700 4865 10734 4899
rect 10768 4865 10802 4899
rect 10836 4865 10870 4899
rect 10904 4865 10938 4899
rect 10972 4865 11006 4899
rect 11040 4865 11074 4899
rect 11108 4865 11142 4899
rect 11176 4865 11210 4899
rect 11244 4865 11278 4899
rect 11312 4865 11346 4899
rect 11380 4865 11414 4899
rect 11448 4865 11482 4899
rect 11516 4865 11550 4899
rect 11584 4865 11618 4899
rect 11652 4865 11686 4899
rect 11720 4865 11754 4899
rect 11788 4865 11822 4899
rect 11856 4865 11890 4899
rect 11924 4865 12071 4899
rect -17 4776 17 4858
rect 51 4824 161 4858
rect 195 4824 229 4858
rect 263 4824 297 4858
rect 331 4824 365 4858
rect 399 4824 433 4858
rect 467 4824 501 4858
rect 535 4824 569 4858
rect 603 4824 637 4858
rect 671 4824 705 4858
rect 739 4824 773 4858
rect 807 4824 841 4858
rect 875 4824 909 4858
rect 943 4824 977 4858
rect 1011 4824 1045 4858
rect 1079 4824 1113 4858
rect 1147 4824 1181 4858
rect 1215 4824 1249 4858
rect 1283 4824 1317 4858
rect 1351 4824 1385 4858
rect 1419 4824 1453 4858
rect 1487 4824 1521 4858
rect 1555 4824 1589 4858
rect 1623 4824 1657 4858
rect 1691 4824 1725 4858
rect 1759 4824 1793 4858
rect 1827 4824 1861 4858
rect 1895 4824 1929 4858
rect 1963 4824 1997 4858
rect 2031 4824 2065 4858
rect 2099 4824 2133 4858
rect 2167 4824 2201 4858
rect 2235 4824 2269 4858
rect 2303 4824 2337 4858
rect 2371 4824 2405 4858
rect 2439 4824 2473 4858
rect 2507 4824 2541 4858
rect 2575 4824 2609 4858
rect 2643 4824 2677 4858
rect 2711 4824 2745 4858
rect 2779 4824 2813 4858
rect 2847 4824 2881 4858
rect 2915 4824 2949 4858
rect 2983 4824 3017 4858
rect 3051 4824 3085 4858
rect 3119 4824 3153 4858
rect 3187 4824 3221 4858
rect 3255 4824 3289 4858
rect 3323 4824 3357 4858
rect 3391 4824 3425 4858
rect 3459 4824 3493 4858
rect 3527 4824 3561 4858
rect 3595 4824 3629 4858
rect 3663 4824 3697 4858
rect 3731 4824 3765 4858
rect 3799 4824 3833 4858
rect 3867 4824 3901 4858
rect 3935 4824 3969 4858
rect 4003 4824 4037 4858
rect 4071 4824 4105 4858
rect 4139 4824 4173 4858
rect 4207 4824 4241 4858
rect 4275 4824 4309 4858
rect 4343 4824 4377 4858
rect 4411 4824 4445 4858
rect 4479 4824 4513 4858
rect 4547 4824 4581 4858
rect 4615 4824 4649 4858
rect 4683 4824 4717 4858
rect 4751 4824 4785 4858
rect 4819 4824 4853 4858
rect 4887 4824 4921 4858
rect 4955 4824 4989 4858
rect 5023 4824 5057 4858
rect 5091 4824 5125 4858
rect 5159 4824 5193 4858
rect 5227 4824 5261 4858
rect 5295 4824 5329 4858
rect 5363 4824 5397 4858
rect 5431 4824 5465 4858
rect 5499 4824 5533 4858
rect 5567 4824 5601 4858
rect 5635 4824 5669 4858
rect 5703 4824 5737 4858
rect 5771 4824 5805 4858
rect 5839 4824 5873 4858
rect 5907 4824 5941 4858
rect 5975 4824 6009 4858
rect 6043 4824 6077 4858
rect 6111 4824 6145 4858
rect 6179 4824 6213 4858
rect 6247 4824 6281 4858
rect 6315 4824 6349 4858
rect 6383 4824 6417 4858
rect 6451 4824 6485 4858
rect 6519 4824 6553 4858
rect 6587 4824 6621 4858
rect 6655 4824 6689 4858
rect 6723 4824 6757 4858
rect 6791 4824 6825 4858
rect 6859 4824 6893 4858
rect 6927 4824 6961 4858
rect 6995 4824 7029 4858
rect 7063 4824 7097 4858
rect 7131 4824 7165 4858
rect 7199 4824 7233 4858
rect 7267 4824 7301 4858
rect 7335 4824 7369 4858
rect 7403 4824 7437 4858
rect 7471 4824 7505 4858
rect 7539 4824 7573 4858
rect 7607 4824 7641 4858
rect 7675 4824 7709 4858
rect 7743 4824 7810 4858
rect -17 4708 17 4742
rect -17 4640 17 4674
rect -17 4572 17 4606
rect 12105 4784 12139 4899
rect 12105 4716 12139 4750
rect 12105 4648 12139 4682
rect -17 4504 17 4538
rect -17 4436 17 4470
rect 321 4411 345 4581
rect 787 4411 811 4581
rect 12105 4580 12139 4614
rect 12105 4512 12139 4546
rect 12078 4444 12139 4478
rect 12078 4417 12112 4444
rect -17 4368 17 4402
rect -17 4300 17 4334
rect -17 4232 17 4266
rect -17 4164 17 4198
rect -17 4096 17 4130
rect -17 4028 17 4062
rect -17 3960 17 3994
rect -17 3892 17 3926
rect -17 3824 17 3858
rect -17 3756 17 3790
rect -17 3688 17 3722
rect -17 3620 17 3654
rect -17 3552 17 3586
rect -17 3484 17 3518
rect 12078 4349 12112 4383
rect 12078 4281 12112 4315
rect 12078 4213 12112 4247
rect 12078 4145 12112 4179
rect 12078 4077 12112 4111
rect 12078 4009 12112 4043
rect 12078 3941 12112 3975
rect 12078 3873 12112 3907
rect 12078 3805 12112 3839
rect 12078 3737 12112 3771
rect 12078 3669 12112 3703
rect 12078 3601 12112 3635
rect 12078 3533 12112 3567
rect -17 3416 17 3450
rect -17 3348 17 3382
rect -17 3280 17 3314
rect -17 3212 17 3246
rect -17 3144 17 3178
rect -17 3076 17 3110
rect -17 3008 17 3042
rect -17 2940 17 2974
rect -17 2872 17 2906
rect 12078 3465 12112 3499
rect 12078 3397 12112 3431
rect 12078 3329 12112 3363
rect 12078 3261 12112 3295
rect 12078 3193 12112 3227
rect 12078 3125 12112 3159
rect 12078 3057 12112 3091
rect 12078 2989 12112 3023
rect 12078 2921 12112 2955
rect -17 2804 17 2838
rect -17 2736 17 2770
rect -17 2668 17 2702
rect -17 2600 17 2634
rect -17 2532 17 2566
rect -17 2464 17 2498
rect -17 2396 17 2430
rect -17 2328 17 2362
rect -17 2260 17 2294
rect 12078 2853 12112 2887
rect 12078 2785 12112 2819
rect 12078 2717 12112 2751
rect 12078 2649 12112 2683
rect 12078 2581 12112 2615
rect 12078 2513 12112 2547
rect 12078 2445 12112 2479
rect 12078 2377 12112 2411
rect 12078 2309 12112 2343
rect -17 2192 17 2226
rect 10154 2245 10188 2269
rect -17 2124 17 2158
rect 3176 2174 4464 2182
rect 3176 2140 3200 2174
rect 3234 2140 3271 2174
rect 3305 2140 3342 2174
rect 3376 2140 3413 2174
rect 3447 2140 3484 2174
rect 3518 2140 3555 2174
rect 3589 2140 3626 2174
rect 3660 2140 3697 2174
rect 3731 2140 3768 2174
rect 3802 2140 3839 2174
rect 3873 2140 3910 2174
rect 3944 2140 3981 2174
rect 4015 2140 4052 2174
rect 4086 2140 4123 2174
rect 4157 2140 4194 2174
rect 4228 2140 4265 2174
rect 4299 2140 4336 2174
rect 4370 2140 4406 2174
rect 4440 2140 4464 2174
rect 3176 2132 4464 2140
rect 10154 2177 10188 2211
rect -17 2056 17 2090
rect -17 1988 17 2022
rect 10154 2109 10188 2143
rect 10154 2041 10188 2075
rect 10154 1973 10188 2007
rect -17 1920 17 1954
rect -17 1852 17 1886
rect -17 1784 17 1818
rect -17 1716 17 1750
rect -17 1648 17 1682
rect -17 1580 17 1614
rect -17 1512 17 1546
rect -17 1444 17 1478
rect -17 1376 17 1410
rect -17 1308 17 1342
rect -17 1240 17 1274
rect -17 1172 17 1206
rect -17 1104 17 1138
rect -17 1036 17 1070
rect 9155 1930 9221 1954
rect 9155 1896 9171 1930
rect 9205 1896 9221 1930
rect 9155 1829 9221 1896
rect 9155 1795 9171 1829
rect 9205 1795 9221 1829
rect 9155 1728 9221 1795
rect 10154 1905 10188 1939
rect 10154 1837 10188 1871
rect 10154 1779 10188 1803
rect 12078 2241 12112 2275
rect 12078 2173 12112 2207
rect 12078 2105 12112 2139
rect 12078 2037 12112 2071
rect 12078 1969 12112 2003
rect 12078 1901 12112 1935
rect 12078 1833 12112 1867
rect 9155 1694 9171 1728
rect 9205 1694 9221 1728
rect 9155 1670 9221 1694
rect 12078 1765 12112 1799
rect 12078 1697 12112 1731
rect 12078 1629 12112 1663
rect 12078 1561 12112 1595
rect 12078 1493 12112 1527
rect 12078 1425 12112 1459
rect 12078 1357 12112 1391
rect 12078 1289 12112 1323
rect 12078 1221 12112 1255
rect 12078 1153 12112 1187
rect 12078 1085 12112 1119
rect -17 968 17 1002
rect -17 900 17 934
rect -17 832 17 866
rect 12078 1017 12112 1051
rect 12078 949 12112 983
rect 12078 881 12112 915
rect 17 810 10605 814
rect 17 798 10472 810
rect -17 781 10472 798
rect -17 747 121 781
rect 155 747 189 781
rect 223 747 257 781
rect 291 747 325 781
rect 359 747 393 781
rect 427 747 461 781
rect 495 747 529 781
rect 563 747 597 781
rect 631 747 665 781
rect 699 747 733 781
rect 767 747 801 781
rect 835 747 869 781
rect 903 747 937 781
rect 971 747 1005 781
rect 1039 747 1073 781
rect 1107 747 1141 781
rect 1175 747 1209 781
rect 1243 747 1277 781
rect 1311 747 1345 781
rect 1379 747 1413 781
rect 1447 747 1481 781
rect 1515 747 1549 781
rect 1583 747 1617 781
rect 1651 747 1685 781
rect 1719 747 1753 781
rect 1787 747 1821 781
rect 1855 747 1889 781
rect 1923 747 1957 781
rect 1991 747 2025 781
rect 2059 747 2093 781
rect 2127 747 2161 781
rect 2195 747 2229 781
rect 2263 747 2297 781
rect 2331 747 2365 781
rect 2399 747 2433 781
rect 2467 747 2501 781
rect 2535 747 2569 781
rect 2603 747 2637 781
rect 2671 747 2705 781
rect 2739 747 2773 781
rect 2807 747 2841 781
rect 2875 747 2909 781
rect 2943 747 2977 781
rect 3011 747 3045 781
rect 3079 747 3113 781
rect 3147 747 3181 781
rect 3215 747 3249 781
rect 3283 747 3317 781
rect 3351 747 3385 781
rect 3419 747 3453 781
rect 3487 747 3521 781
rect 3555 747 3589 781
rect 3623 747 3657 781
rect 3691 747 3725 781
rect 3759 747 3793 781
rect 3827 747 3861 781
rect 3895 747 3929 781
rect 3963 747 3997 781
rect 4031 747 4065 781
rect 4099 747 4133 781
rect 4167 747 4201 781
rect 4235 747 4269 781
rect 4303 747 4337 781
rect 4371 747 4405 781
rect 4439 747 4473 781
rect 4507 747 4541 781
rect 4575 747 4609 781
rect 4643 747 4677 781
rect 4711 747 4745 781
rect 4779 747 4813 781
rect 4847 747 4881 781
rect 4915 747 4949 781
rect 4983 747 5017 781
rect 5051 747 5085 781
rect 5119 747 5153 781
rect 5187 747 5221 781
rect 5255 747 5289 781
rect 5323 747 5357 781
rect 5391 747 5425 781
rect 5459 747 5493 781
rect 5527 747 5561 781
rect 5595 747 5629 781
rect 5663 747 5697 781
rect 5731 747 5765 781
rect 5799 747 5833 781
rect 5867 747 5901 781
rect 5935 747 5969 781
rect 6003 747 6037 781
rect 6071 747 6105 781
rect 6139 747 6173 781
rect 6207 747 6241 781
rect 6275 747 6309 781
rect 6343 747 6377 781
rect 6411 747 6445 781
rect 6479 747 6513 781
rect 6547 747 6581 781
rect 6615 747 6649 781
rect 6683 747 6717 781
rect 6751 747 6785 781
rect 6819 747 6853 781
rect 6887 747 6921 781
rect 6955 747 6989 781
rect 7023 747 7057 781
rect 7091 747 7125 781
rect 7159 747 7193 781
rect 7227 747 7261 781
rect 7295 747 7329 781
rect 7363 747 7397 781
rect 7431 747 7465 781
rect 7499 747 7533 781
rect 7567 747 7601 781
rect 7635 747 7669 781
rect 7703 747 7737 781
rect 7771 747 7805 781
rect 7839 747 7873 781
rect 7907 747 7941 781
rect 7975 747 8009 781
rect 8043 747 8077 781
rect 8111 747 8145 781
rect 8179 747 8213 781
rect 8247 747 8281 781
rect 8315 747 8349 781
rect 8383 747 8417 781
rect 8451 747 8485 781
rect 8519 747 8553 781
rect 8587 747 8621 781
rect 8655 747 8689 781
rect 8723 747 8757 781
rect 8791 747 8825 781
rect 8859 747 8893 781
rect 8927 747 8961 781
rect 8995 747 9029 781
rect 9063 747 9097 781
rect 9131 747 9165 781
rect 9199 747 9233 781
rect 9267 747 9301 781
rect 9335 747 9369 781
rect 9403 747 9437 781
rect 9471 747 9505 781
rect 9539 747 9573 781
rect 9607 747 9641 781
rect 9675 747 9709 781
rect 9743 747 9777 781
rect 9811 747 9845 781
rect 9879 747 9913 781
rect 9947 747 9981 781
rect 10015 747 10049 781
rect 10083 747 10117 781
rect 10151 747 10185 781
rect 10219 747 10253 781
rect 10287 747 10321 781
rect 10355 776 10472 781
rect 10506 776 10605 810
rect 10355 747 10605 776
rect -17 735 10605 747
rect -17 714 10551 735
rect 10505 701 10551 714
rect 10585 701 10605 735
rect 10505 677 10605 701
rect 12078 813 12112 847
rect 12078 745 12112 779
rect 12078 677 12112 711
rect 10505 661 12112 677
rect 10505 627 10621 661
rect 10655 627 10692 661
rect 10726 627 10763 661
rect 10797 627 10834 661
rect 10868 627 10905 661
rect 10939 627 10976 661
rect 11010 627 11047 661
rect 11081 627 11118 661
rect 11152 627 11189 661
rect 11223 627 11260 661
rect 11294 627 11331 661
rect 11365 627 11402 661
rect 11436 627 11473 661
rect 11507 627 11544 661
rect 11578 627 11615 661
rect 11649 627 11686 661
rect 11720 627 11757 661
rect 11791 627 11828 661
rect 11862 627 11899 661
rect 11933 627 11970 661
rect 12004 627 12041 661
rect 12075 627 12112 661
rect 10505 565 12112 627
<< mvpsubdiffcont >>
rect 9157 3441 9191 3475
rect 9225 3441 9259 3475
rect 9157 3367 9191 3401
rect 9225 3367 9259 3401
rect 9157 3293 9191 3327
rect 9225 3293 9259 3327
rect 9157 3219 9191 3253
rect 9225 3219 9259 3253
rect 9157 3145 9191 3179
rect 9225 3145 9259 3179
rect 9157 3071 9191 3105
rect 9225 3071 9259 3105
rect 9157 2997 9191 3031
rect 9225 2997 9259 3031
rect 9157 2923 9191 2957
rect 9225 2923 9259 2957
rect 8463 1896 8497 1930
rect 8563 1896 8597 1930
rect 8663 1896 8697 1930
rect 8463 1822 8497 1856
rect 8563 1822 8597 1856
rect 8663 1822 8697 1856
rect 8463 1748 8497 1782
rect 8563 1748 8597 1782
rect 8663 1748 8697 1782
rect 8463 1674 8497 1708
rect 8563 1674 8597 1708
rect 8663 1674 8697 1708
rect 8463 1600 8497 1634
rect 8563 1600 8597 1634
rect 8663 1600 8697 1634
rect 8463 1526 8497 1560
rect 8563 1526 8597 1560
rect 8663 1526 8697 1560
rect 8463 1453 8497 1487
rect 8563 1453 8597 1487
rect 8663 1453 8697 1487
rect 8463 1380 8497 1414
rect 8563 1380 8597 1414
rect 8663 1380 8697 1414
rect 8463 1307 8497 1341
rect 8563 1307 8597 1341
rect 8663 1307 8697 1341
rect 8463 1234 8497 1268
rect 8563 1234 8597 1268
rect 8663 1234 8697 1268
rect 8463 1161 8497 1195
rect 8563 1161 8597 1195
rect 8663 1161 8697 1195
rect 8463 1088 8497 1122
rect 8563 1088 8597 1122
rect 8663 1088 8697 1122
<< mvnsubdiffcont >>
rect 7810 4865 7844 4899
rect 7878 4865 7912 4899
rect 7946 4865 7980 4899
rect 8014 4865 8048 4899
rect 8082 4865 8116 4899
rect 8150 4865 8184 4899
rect 8218 4865 8252 4899
rect 8286 4865 8320 4899
rect 8354 4865 8388 4899
rect 8422 4865 8456 4899
rect 8490 4865 8524 4899
rect 8558 4865 8592 4899
rect 8626 4865 8660 4899
rect 8694 4865 8728 4899
rect 8762 4865 8796 4899
rect 8830 4865 8864 4899
rect 8898 4865 8932 4899
rect 8966 4865 9000 4899
rect 9034 4865 9068 4899
rect 9102 4865 9136 4899
rect 9170 4865 9204 4899
rect 9238 4865 9272 4899
rect 9306 4865 9340 4899
rect 9374 4865 9408 4899
rect 9442 4865 9476 4899
rect 9510 4865 9544 4899
rect 9578 4865 9612 4899
rect 9646 4865 9680 4899
rect 9714 4865 9748 4899
rect 9782 4865 9816 4899
rect 9850 4865 9884 4899
rect 9918 4865 9952 4899
rect 9986 4865 10020 4899
rect 10054 4865 10088 4899
rect 10122 4865 10156 4899
rect 10190 4865 10224 4899
rect 10258 4865 10292 4899
rect 10326 4865 10360 4899
rect 10394 4865 10428 4899
rect 10462 4865 10496 4899
rect 10530 4865 10564 4899
rect 10598 4865 10632 4899
rect 10666 4865 10700 4899
rect 10734 4865 10768 4899
rect 10802 4865 10836 4899
rect 10870 4865 10904 4899
rect 10938 4865 10972 4899
rect 11006 4865 11040 4899
rect 11074 4865 11108 4899
rect 11142 4865 11176 4899
rect 11210 4865 11244 4899
rect 11278 4865 11312 4899
rect 11346 4865 11380 4899
rect 11414 4865 11448 4899
rect 11482 4865 11516 4899
rect 11550 4865 11584 4899
rect 11618 4865 11652 4899
rect 11686 4865 11720 4899
rect 11754 4865 11788 4899
rect 11822 4865 11856 4899
rect 11890 4865 11924 4899
rect 12071 4865 12105 4899
rect 17 4824 51 4858
rect 161 4824 195 4858
rect 229 4824 263 4858
rect 297 4824 331 4858
rect 365 4824 399 4858
rect 433 4824 467 4858
rect 501 4824 535 4858
rect 569 4824 603 4858
rect 637 4824 671 4858
rect 705 4824 739 4858
rect 773 4824 807 4858
rect 841 4824 875 4858
rect 909 4824 943 4858
rect 977 4824 1011 4858
rect 1045 4824 1079 4858
rect 1113 4824 1147 4858
rect 1181 4824 1215 4858
rect 1249 4824 1283 4858
rect 1317 4824 1351 4858
rect 1385 4824 1419 4858
rect 1453 4824 1487 4858
rect 1521 4824 1555 4858
rect 1589 4824 1623 4858
rect 1657 4824 1691 4858
rect 1725 4824 1759 4858
rect 1793 4824 1827 4858
rect 1861 4824 1895 4858
rect 1929 4824 1963 4858
rect 1997 4824 2031 4858
rect 2065 4824 2099 4858
rect 2133 4824 2167 4858
rect 2201 4824 2235 4858
rect 2269 4824 2303 4858
rect 2337 4824 2371 4858
rect 2405 4824 2439 4858
rect 2473 4824 2507 4858
rect 2541 4824 2575 4858
rect 2609 4824 2643 4858
rect 2677 4824 2711 4858
rect 2745 4824 2779 4858
rect 2813 4824 2847 4858
rect 2881 4824 2915 4858
rect 2949 4824 2983 4858
rect 3017 4824 3051 4858
rect 3085 4824 3119 4858
rect 3153 4824 3187 4858
rect 3221 4824 3255 4858
rect 3289 4824 3323 4858
rect 3357 4824 3391 4858
rect 3425 4824 3459 4858
rect 3493 4824 3527 4858
rect 3561 4824 3595 4858
rect 3629 4824 3663 4858
rect 3697 4824 3731 4858
rect 3765 4824 3799 4858
rect 3833 4824 3867 4858
rect 3901 4824 3935 4858
rect 3969 4824 4003 4858
rect 4037 4824 4071 4858
rect 4105 4824 4139 4858
rect 4173 4824 4207 4858
rect 4241 4824 4275 4858
rect 4309 4824 4343 4858
rect 4377 4824 4411 4858
rect 4445 4824 4479 4858
rect 4513 4824 4547 4858
rect 4581 4824 4615 4858
rect 4649 4824 4683 4858
rect 4717 4824 4751 4858
rect 4785 4824 4819 4858
rect 4853 4824 4887 4858
rect 4921 4824 4955 4858
rect 4989 4824 5023 4858
rect 5057 4824 5091 4858
rect 5125 4824 5159 4858
rect 5193 4824 5227 4858
rect 5261 4824 5295 4858
rect 5329 4824 5363 4858
rect 5397 4824 5431 4858
rect 5465 4824 5499 4858
rect 5533 4824 5567 4858
rect 5601 4824 5635 4858
rect 5669 4824 5703 4858
rect 5737 4824 5771 4858
rect 5805 4824 5839 4858
rect 5873 4824 5907 4858
rect 5941 4824 5975 4858
rect 6009 4824 6043 4858
rect 6077 4824 6111 4858
rect 6145 4824 6179 4858
rect 6213 4824 6247 4858
rect 6281 4824 6315 4858
rect 6349 4824 6383 4858
rect 6417 4824 6451 4858
rect 6485 4824 6519 4858
rect 6553 4824 6587 4858
rect 6621 4824 6655 4858
rect 6689 4824 6723 4858
rect 6757 4824 6791 4858
rect 6825 4824 6859 4858
rect 6893 4824 6927 4858
rect 6961 4824 6995 4858
rect 7029 4824 7063 4858
rect 7097 4824 7131 4858
rect 7165 4824 7199 4858
rect 7233 4824 7267 4858
rect 7301 4824 7335 4858
rect 7369 4824 7403 4858
rect 7437 4824 7471 4858
rect 7505 4824 7539 4858
rect 7573 4824 7607 4858
rect 7641 4824 7675 4858
rect 7709 4824 7743 4858
rect -17 4742 17 4776
rect -17 4674 17 4708
rect -17 4606 17 4640
rect 12105 4750 12139 4784
rect 12105 4682 12139 4716
rect 12105 4614 12139 4648
rect -17 4538 17 4572
rect -17 4470 17 4504
rect -17 4402 17 4436
rect 345 4411 787 4581
rect 12105 4546 12139 4580
rect 12105 4478 12139 4512
rect -17 4334 17 4368
rect -17 4266 17 4300
rect -17 4198 17 4232
rect -17 4130 17 4164
rect -17 4062 17 4096
rect -17 3994 17 4028
rect -17 3926 17 3960
rect -17 3858 17 3892
rect -17 3790 17 3824
rect -17 3722 17 3756
rect -17 3654 17 3688
rect -17 3586 17 3620
rect -17 3518 17 3552
rect 12078 4383 12112 4417
rect 12078 4315 12112 4349
rect 12078 4247 12112 4281
rect 12078 4179 12112 4213
rect 12078 4111 12112 4145
rect 12078 4043 12112 4077
rect 12078 3975 12112 4009
rect 12078 3907 12112 3941
rect 12078 3839 12112 3873
rect 12078 3771 12112 3805
rect 12078 3703 12112 3737
rect 12078 3635 12112 3669
rect 12078 3567 12112 3601
rect 12078 3499 12112 3533
rect -17 3450 17 3484
rect -17 3382 17 3416
rect -17 3314 17 3348
rect -17 3246 17 3280
rect -17 3178 17 3212
rect -17 3110 17 3144
rect -17 3042 17 3076
rect -17 2974 17 3008
rect -17 2906 17 2940
rect 12078 3431 12112 3465
rect 12078 3363 12112 3397
rect 12078 3295 12112 3329
rect 12078 3227 12112 3261
rect 12078 3159 12112 3193
rect 12078 3091 12112 3125
rect 12078 3023 12112 3057
rect 12078 2955 12112 2989
rect -17 2838 17 2872
rect -17 2770 17 2804
rect -17 2702 17 2736
rect -17 2634 17 2668
rect -17 2566 17 2600
rect -17 2498 17 2532
rect -17 2430 17 2464
rect -17 2362 17 2396
rect -17 2294 17 2328
rect 12078 2887 12112 2921
rect 12078 2819 12112 2853
rect 12078 2751 12112 2785
rect 12078 2683 12112 2717
rect 12078 2615 12112 2649
rect 12078 2547 12112 2581
rect 12078 2479 12112 2513
rect 12078 2411 12112 2445
rect 12078 2343 12112 2377
rect 12078 2275 12112 2309
rect -17 2226 17 2260
rect -17 2158 17 2192
rect 10154 2211 10188 2245
rect 3200 2140 3234 2174
rect 3271 2140 3305 2174
rect 3342 2140 3376 2174
rect 3413 2140 3447 2174
rect 3484 2140 3518 2174
rect 3555 2140 3589 2174
rect 3626 2140 3660 2174
rect 3697 2140 3731 2174
rect 3768 2140 3802 2174
rect 3839 2140 3873 2174
rect 3910 2140 3944 2174
rect 3981 2140 4015 2174
rect 4052 2140 4086 2174
rect 4123 2140 4157 2174
rect 4194 2140 4228 2174
rect 4265 2140 4299 2174
rect 4336 2140 4370 2174
rect 4406 2140 4440 2174
rect 10154 2143 10188 2177
rect -17 2090 17 2124
rect -17 2022 17 2056
rect -17 1954 17 1988
rect 10154 2075 10188 2109
rect 10154 2007 10188 2041
rect -17 1886 17 1920
rect -17 1818 17 1852
rect -17 1750 17 1784
rect -17 1682 17 1716
rect -17 1614 17 1648
rect -17 1546 17 1580
rect -17 1478 17 1512
rect -17 1410 17 1444
rect -17 1342 17 1376
rect -17 1274 17 1308
rect -17 1206 17 1240
rect -17 1138 17 1172
rect -17 1070 17 1104
rect 9171 1896 9205 1930
rect 9171 1795 9205 1829
rect 10154 1939 10188 1973
rect 10154 1871 10188 1905
rect 10154 1803 10188 1837
rect 12078 2207 12112 2241
rect 12078 2139 12112 2173
rect 12078 2071 12112 2105
rect 12078 2003 12112 2037
rect 12078 1935 12112 1969
rect 12078 1867 12112 1901
rect 12078 1799 12112 1833
rect 9171 1694 9205 1728
rect 12078 1731 12112 1765
rect 12078 1663 12112 1697
rect 12078 1595 12112 1629
rect 12078 1527 12112 1561
rect 12078 1459 12112 1493
rect 12078 1391 12112 1425
rect 12078 1323 12112 1357
rect 12078 1255 12112 1289
rect 12078 1187 12112 1221
rect 12078 1119 12112 1153
rect -17 1002 17 1036
rect -17 934 17 968
rect -17 866 17 900
rect -17 798 17 832
rect 12078 1051 12112 1085
rect 12078 983 12112 1017
rect 12078 915 12112 949
rect 12078 847 12112 881
rect 121 747 155 781
rect 189 747 223 781
rect 257 747 291 781
rect 325 747 359 781
rect 393 747 427 781
rect 461 747 495 781
rect 529 747 563 781
rect 597 747 631 781
rect 665 747 699 781
rect 733 747 767 781
rect 801 747 835 781
rect 869 747 903 781
rect 937 747 971 781
rect 1005 747 1039 781
rect 1073 747 1107 781
rect 1141 747 1175 781
rect 1209 747 1243 781
rect 1277 747 1311 781
rect 1345 747 1379 781
rect 1413 747 1447 781
rect 1481 747 1515 781
rect 1549 747 1583 781
rect 1617 747 1651 781
rect 1685 747 1719 781
rect 1753 747 1787 781
rect 1821 747 1855 781
rect 1889 747 1923 781
rect 1957 747 1991 781
rect 2025 747 2059 781
rect 2093 747 2127 781
rect 2161 747 2195 781
rect 2229 747 2263 781
rect 2297 747 2331 781
rect 2365 747 2399 781
rect 2433 747 2467 781
rect 2501 747 2535 781
rect 2569 747 2603 781
rect 2637 747 2671 781
rect 2705 747 2739 781
rect 2773 747 2807 781
rect 2841 747 2875 781
rect 2909 747 2943 781
rect 2977 747 3011 781
rect 3045 747 3079 781
rect 3113 747 3147 781
rect 3181 747 3215 781
rect 3249 747 3283 781
rect 3317 747 3351 781
rect 3385 747 3419 781
rect 3453 747 3487 781
rect 3521 747 3555 781
rect 3589 747 3623 781
rect 3657 747 3691 781
rect 3725 747 3759 781
rect 3793 747 3827 781
rect 3861 747 3895 781
rect 3929 747 3963 781
rect 3997 747 4031 781
rect 4065 747 4099 781
rect 4133 747 4167 781
rect 4201 747 4235 781
rect 4269 747 4303 781
rect 4337 747 4371 781
rect 4405 747 4439 781
rect 4473 747 4507 781
rect 4541 747 4575 781
rect 4609 747 4643 781
rect 4677 747 4711 781
rect 4745 747 4779 781
rect 4813 747 4847 781
rect 4881 747 4915 781
rect 4949 747 4983 781
rect 5017 747 5051 781
rect 5085 747 5119 781
rect 5153 747 5187 781
rect 5221 747 5255 781
rect 5289 747 5323 781
rect 5357 747 5391 781
rect 5425 747 5459 781
rect 5493 747 5527 781
rect 5561 747 5595 781
rect 5629 747 5663 781
rect 5697 747 5731 781
rect 5765 747 5799 781
rect 5833 747 5867 781
rect 5901 747 5935 781
rect 5969 747 6003 781
rect 6037 747 6071 781
rect 6105 747 6139 781
rect 6173 747 6207 781
rect 6241 747 6275 781
rect 6309 747 6343 781
rect 6377 747 6411 781
rect 6445 747 6479 781
rect 6513 747 6547 781
rect 6581 747 6615 781
rect 6649 747 6683 781
rect 6717 747 6751 781
rect 6785 747 6819 781
rect 6853 747 6887 781
rect 6921 747 6955 781
rect 6989 747 7023 781
rect 7057 747 7091 781
rect 7125 747 7159 781
rect 7193 747 7227 781
rect 7261 747 7295 781
rect 7329 747 7363 781
rect 7397 747 7431 781
rect 7465 747 7499 781
rect 7533 747 7567 781
rect 7601 747 7635 781
rect 7669 747 7703 781
rect 7737 747 7771 781
rect 7805 747 7839 781
rect 7873 747 7907 781
rect 7941 747 7975 781
rect 8009 747 8043 781
rect 8077 747 8111 781
rect 8145 747 8179 781
rect 8213 747 8247 781
rect 8281 747 8315 781
rect 8349 747 8383 781
rect 8417 747 8451 781
rect 8485 747 8519 781
rect 8553 747 8587 781
rect 8621 747 8655 781
rect 8689 747 8723 781
rect 8757 747 8791 781
rect 8825 747 8859 781
rect 8893 747 8927 781
rect 8961 747 8995 781
rect 9029 747 9063 781
rect 9097 747 9131 781
rect 9165 747 9199 781
rect 9233 747 9267 781
rect 9301 747 9335 781
rect 9369 747 9403 781
rect 9437 747 9471 781
rect 9505 747 9539 781
rect 9573 747 9607 781
rect 9641 747 9675 781
rect 9709 747 9743 781
rect 9777 747 9811 781
rect 9845 747 9879 781
rect 9913 747 9947 781
rect 9981 747 10015 781
rect 10049 747 10083 781
rect 10117 747 10151 781
rect 10185 747 10219 781
rect 10253 747 10287 781
rect 10321 747 10355 781
rect 10472 776 10506 810
rect 10551 701 10585 735
rect 12078 779 12112 813
rect 12078 711 12112 745
rect 10621 627 10655 661
rect 10692 627 10726 661
rect 10763 627 10797 661
rect 10834 627 10868 661
rect 10905 627 10939 661
rect 10976 627 11010 661
rect 11047 627 11081 661
rect 11118 627 11152 661
rect 11189 627 11223 661
rect 11260 627 11294 661
rect 11331 627 11365 661
rect 11402 627 11436 661
rect 11473 627 11507 661
rect 11544 627 11578 661
rect 11615 627 11649 661
rect 11686 627 11720 661
rect 11757 627 11791 661
rect 11828 627 11862 661
rect 11899 627 11933 661
rect 11970 627 12004 661
rect 12041 627 12075 661
<< locali >>
rect 7776 4858 7810 4899
rect 7844 4865 7878 4899
rect 7912 4865 7946 4899
rect 7980 4865 8014 4899
rect 8048 4865 8082 4899
rect 8116 4865 8150 4899
rect 8184 4865 8218 4899
rect 8252 4865 8286 4899
rect 8320 4865 8354 4899
rect 8388 4865 8422 4899
rect 8456 4865 8490 4899
rect 8524 4865 8558 4899
rect 8592 4865 8626 4899
rect 8660 4865 8694 4899
rect 8728 4865 8762 4899
rect 8796 4865 8830 4899
rect 8864 4865 8898 4899
rect 8932 4865 8966 4899
rect 9000 4865 9034 4899
rect 9068 4865 9102 4899
rect 9136 4865 9170 4899
rect 9204 4865 9238 4899
rect 9272 4865 9306 4899
rect 9340 4865 9374 4899
rect 9408 4865 9442 4899
rect 9476 4865 9510 4899
rect 9544 4865 9578 4899
rect 9612 4865 9646 4899
rect 9680 4865 9714 4899
rect 9748 4865 9782 4899
rect 9816 4865 9850 4899
rect 9884 4865 9918 4899
rect 9952 4865 9986 4899
rect 10020 4865 10054 4899
rect 10088 4865 10122 4899
rect 10156 4865 10190 4899
rect 10224 4865 10258 4899
rect 10292 4865 10326 4899
rect 10360 4865 10394 4899
rect 10428 4865 10462 4899
rect 10496 4865 10530 4899
rect 10564 4865 10598 4899
rect 10632 4865 10666 4899
rect 10700 4865 10734 4899
rect 10768 4865 10802 4899
rect 10836 4865 10870 4899
rect 10904 4865 10938 4899
rect 10972 4865 11006 4899
rect 11040 4865 11074 4899
rect 11108 4865 11142 4899
rect 11176 4865 11210 4899
rect 11244 4865 11278 4899
rect 11312 4865 11346 4899
rect 11380 4865 11414 4899
rect 11448 4865 11482 4899
rect 11516 4865 11550 4899
rect 11584 4865 11618 4899
rect 11652 4865 11686 4899
rect 11720 4865 11754 4899
rect 11788 4865 11822 4899
rect 11856 4865 11890 4899
rect 11924 4865 12071 4899
rect -17 4776 17 4858
rect 51 4824 161 4858
rect 195 4824 229 4858
rect 263 4824 297 4858
rect 331 4824 365 4858
rect 399 4824 433 4858
rect 467 4824 501 4858
rect 535 4824 569 4858
rect 603 4824 637 4858
rect 671 4824 705 4858
rect 739 4824 773 4858
rect 807 4824 841 4858
rect 875 4824 909 4858
rect 943 4824 977 4858
rect 1011 4824 1045 4858
rect 1079 4824 1113 4858
rect 1147 4824 1181 4858
rect 1215 4824 1249 4858
rect 1283 4824 1317 4858
rect 1351 4824 1385 4858
rect 1419 4824 1453 4858
rect 1487 4824 1521 4858
rect 1555 4824 1589 4858
rect 1623 4824 1657 4858
rect 1691 4824 1725 4858
rect 1759 4824 1793 4858
rect 1827 4824 1861 4858
rect 1895 4824 1929 4858
rect 1963 4824 1997 4858
rect 2031 4824 2065 4858
rect 2099 4824 2133 4858
rect 2167 4824 2201 4858
rect 2235 4824 2269 4858
rect 2303 4824 2337 4858
rect 2371 4824 2405 4858
rect 2439 4824 2473 4858
rect 2507 4824 2541 4858
rect 2575 4824 2609 4858
rect 2643 4824 2677 4858
rect 2711 4824 2745 4858
rect 2779 4824 2813 4858
rect 2847 4824 2881 4858
rect 2915 4824 2949 4858
rect 2983 4824 3017 4858
rect 3051 4824 3085 4858
rect 3119 4824 3153 4858
rect 3187 4824 3221 4858
rect 3255 4824 3289 4858
rect 3323 4824 3357 4858
rect 3391 4824 3425 4858
rect 3459 4824 3493 4858
rect 3527 4824 3561 4858
rect 3595 4824 3629 4858
rect 3663 4824 3697 4858
rect 3731 4824 3765 4858
rect 3799 4824 3833 4858
rect 3867 4824 3901 4858
rect 3935 4824 3969 4858
rect 4003 4824 4037 4858
rect 4071 4824 4105 4858
rect 4139 4824 4173 4858
rect 4207 4824 4241 4858
rect 4275 4824 4309 4858
rect 4343 4824 4377 4858
rect 4411 4824 4445 4858
rect 4479 4824 4513 4858
rect 4547 4824 4581 4858
rect 4615 4824 4649 4858
rect 4683 4824 4717 4858
rect 4751 4824 4785 4858
rect 4819 4824 4853 4858
rect 4887 4824 4921 4858
rect 4955 4824 4989 4858
rect 5023 4824 5057 4858
rect 5091 4824 5125 4858
rect 5159 4824 5193 4858
rect 5227 4824 5261 4858
rect 5295 4824 5329 4858
rect 5363 4824 5397 4858
rect 5431 4824 5465 4858
rect 5499 4824 5533 4858
rect 5567 4824 5601 4858
rect 5635 4824 5669 4858
rect 5703 4824 5737 4858
rect 5771 4824 5805 4858
rect 5839 4824 5873 4858
rect 5907 4824 5941 4858
rect 5975 4824 6009 4858
rect 6043 4824 6077 4858
rect 6111 4824 6145 4858
rect 6179 4824 6213 4858
rect 6247 4824 6281 4858
rect 6315 4824 6349 4858
rect 6383 4824 6417 4858
rect 6451 4824 6485 4858
rect 6519 4824 6553 4858
rect 6587 4824 6621 4858
rect 6655 4824 6689 4858
rect 6723 4824 6757 4858
rect 6791 4824 6825 4858
rect 6859 4824 6893 4858
rect 6927 4824 6961 4858
rect 6995 4824 7029 4858
rect 7063 4824 7097 4858
rect 7131 4824 7165 4858
rect 7199 4824 7233 4858
rect 7267 4824 7301 4858
rect 7335 4824 7369 4858
rect 7403 4824 7437 4858
rect 7471 4824 7505 4858
rect 7539 4824 7573 4858
rect 7607 4824 7641 4858
rect 7675 4824 7709 4858
rect 7743 4824 7810 4858
rect -17 4708 17 4742
rect 12105 4784 12139 4899
rect 12105 4716 12139 4750
rect -17 4640 17 4674
rect -17 4572 17 4606
rect -17 4504 17 4538
rect -17 4436 17 4470
rect 321 4543 345 4581
rect 787 4543 811 4581
rect 321 4437 333 4543
rect 799 4437 811 4543
rect 321 4411 345 4437
rect 787 4411 811 4437
rect -17 4368 17 4402
rect -17 4300 17 4334
rect -17 4232 17 4266
rect -17 4164 17 4198
rect -17 4096 17 4130
rect -17 4028 17 4062
rect -17 3960 17 3994
rect -17 3892 17 3926
rect -17 3824 17 3858
rect -17 3756 17 3790
rect -17 3688 17 3722
rect 7208 3669 7242 4711
rect 12105 4648 12139 4682
rect 12105 4580 12139 4614
rect 12105 4527 12139 4546
rect 12112 4512 12139 4527
rect 12078 4478 12105 4493
rect 12078 4453 12139 4478
rect 12112 4444 12139 4453
rect 12078 4417 12112 4419
rect 12078 4379 12112 4383
rect 8771 4311 8809 4345
rect 12078 4306 12112 4315
rect 12078 4233 12112 4247
rect 12078 4160 12112 4179
rect 12078 4077 12112 4111
rect 12078 4009 12112 4043
rect 12078 3941 12112 3975
rect 12078 3873 12112 3907
rect 12078 3805 12112 3839
rect 12078 3737 12112 3771
rect -17 3620 17 3654
rect 7122 3635 7138 3669
rect 7172 3635 7210 3669
rect 7244 3635 7256 3669
rect 7122 3605 7256 3635
rect -17 3552 17 3586
rect 7163 3529 7228 3571
rect 7538 3561 7552 3567
rect 7586 3561 7624 3595
rect 7885 3580 7896 3595
rect 7658 3561 7672 3567
rect 7930 3561 7968 3595
rect 8002 3580 8019 3595
rect -17 3484 17 3518
rect -17 3416 17 3450
rect -17 3348 17 3382
rect -17 3280 17 3314
rect -17 3212 17 3246
rect -17 3144 17 3178
rect -17 3076 17 3110
rect -17 3008 17 3042
rect -17 2940 17 2974
rect -17 2872 17 2906
rect -17 2804 17 2838
rect 7164 2861 7228 3529
rect 8183 3521 8385 3556
rect 8183 3487 8259 3521
rect 8293 3487 8331 3521
rect 8365 3487 8385 3521
rect 8648 3519 8831 3548
rect 8648 3485 8659 3519
rect 8693 3485 8731 3519
rect 8765 3485 8831 3519
rect 8884 3504 9067 3691
rect 12078 3669 12112 3703
rect 9440 3642 9454 3669
rect 9434 3635 9454 3642
rect 9488 3635 9526 3669
rect 9560 3635 9598 3669
rect 9632 3635 9670 3669
rect 9132 3580 9144 3595
rect 9178 3561 9216 3595
rect 9250 3580 9266 3595
rect 9434 3582 9704 3635
rect 12078 3601 12112 3635
rect 10031 3549 10069 3583
rect 10103 3549 10141 3583
rect 12078 3533 12112 3567
rect 7164 2817 7449 2861
rect 8757 2851 8831 3485
rect 8899 2895 8970 3476
rect 9157 3475 9259 3499
rect 9191 3441 9225 3475
rect 9157 3401 9259 3441
rect 9191 3372 9225 3401
rect 12078 3465 12112 3499
rect 12078 3397 12112 3431
rect 9157 3179 9259 3194
rect 11792 3333 11814 3367
rect 11848 3333 11870 3367
rect 11792 3295 11870 3333
rect 11792 3261 11814 3295
rect 11848 3261 11870 3295
rect 11792 3223 11870 3261
rect 11792 3189 11814 3223
rect 11848 3189 11870 3223
rect 12078 3360 12112 3363
rect 12078 3284 12112 3295
rect 12078 3208 12112 3227
rect 9191 3145 9225 3179
rect 9157 3105 9259 3145
rect 9191 3071 9225 3105
rect 9157 3031 9259 3071
rect 9191 2997 9225 3031
rect 9157 2957 9259 2997
rect 9191 2923 9225 2957
rect 9157 2899 9259 2923
rect 12078 3132 12112 3159
rect 12078 3057 12112 3091
rect 12078 2989 12112 3022
rect 12078 2921 12112 2946
rect 12078 2853 12112 2870
rect -17 2736 17 2770
rect -17 2668 17 2702
rect -17 2600 17 2634
rect -17 2532 17 2566
rect -17 2464 17 2498
rect -17 2396 17 2430
rect -17 2328 17 2362
rect 12078 2785 12112 2794
rect 12078 2717 12112 2751
rect 12078 2649 12112 2683
rect 12078 2581 12112 2615
rect 12078 2513 12112 2547
rect 12078 2445 12112 2465
rect 12078 2377 12112 2393
rect -17 2260 17 2294
rect 1463 2267 4620 2336
rect 12078 2309 12112 2321
rect 1463 2264 3070 2267
rect 3025 2233 3070 2264
rect 3104 2233 3144 2267
rect 3178 2233 3218 2267
rect 3252 2233 3292 2267
rect 3326 2233 3366 2267
rect 3400 2233 3440 2267
rect 3474 2233 3514 2267
rect 3548 2233 3588 2267
rect 3622 2233 3662 2267
rect 3696 2233 3736 2267
rect 3770 2233 3810 2267
rect 3844 2233 3884 2267
rect 3918 2233 3958 2267
rect 3992 2233 4032 2267
rect 4066 2233 4106 2267
rect 4140 2233 4180 2267
rect 4214 2233 4253 2267
rect 4287 2233 4326 2267
rect 4360 2233 4399 2267
rect 4433 2233 4472 2267
rect 4506 2233 4545 2267
rect 4579 2233 4618 2267
rect 10154 2245 10229 2269
rect -17 2192 17 2226
rect 10188 2211 10229 2245
rect -17 2124 17 2158
rect 3176 2174 4464 2182
rect 3176 2140 3200 2174
rect 3234 2140 3271 2174
rect 3305 2140 3342 2174
rect 3376 2140 3413 2174
rect 3447 2140 3484 2174
rect 3518 2140 3555 2174
rect 3589 2140 3626 2174
rect 3660 2140 3697 2174
rect 3731 2140 3768 2174
rect 3802 2140 3839 2174
rect 3873 2140 3910 2174
rect 3944 2140 3981 2174
rect 4015 2140 4052 2174
rect 4086 2140 4123 2174
rect 4157 2140 4194 2174
rect 4228 2140 4265 2174
rect 4299 2140 4336 2174
rect 4370 2140 4406 2174
rect 4440 2140 4464 2174
rect 3176 2132 4464 2140
rect 10154 2177 10229 2211
rect 10188 2143 10229 2177
rect -17 2056 17 2090
rect -17 1988 17 2022
rect 3316 2008 3350 2132
rect 3628 2008 3662 2132
rect -17 1920 17 1954
rect -17 1852 17 1886
rect -17 1784 17 1818
rect -17 1716 17 1750
rect -17 1648 17 1682
rect -17 1580 17 1614
rect -17 1512 17 1546
rect -17 1444 17 1478
rect -17 1376 17 1410
rect -17 1308 17 1342
rect -17 1240 17 1274
rect -17 1172 17 1206
rect -17 1104 17 1138
rect -17 1036 17 1070
rect 3940 1008 4072 2132
rect 10154 2109 10229 2143
rect 10188 2075 10229 2109
rect 10154 2041 10229 2075
rect 10188 2007 10229 2041
rect 10154 1973 10229 2007
rect 8463 1930 8697 1954
rect 8497 1896 8563 1930
rect 8597 1896 8663 1930
rect 8463 1856 8697 1896
rect 8497 1822 8563 1856
rect 8597 1822 8663 1856
rect 8463 1782 8697 1822
rect 8497 1748 8563 1782
rect 8597 1748 8663 1782
rect 8463 1708 8697 1748
rect 8497 1674 8563 1708
rect 8597 1674 8663 1708
rect 8463 1634 8697 1674
rect 9155 1930 9221 1954
rect 9155 1896 9171 1930
rect 9205 1896 9221 1930
rect 9155 1829 9221 1896
rect 9155 1795 9171 1829
rect 9205 1795 9221 1829
rect 9155 1728 9221 1795
rect 10188 1939 10229 1973
rect 10154 1905 10229 1939
rect 10188 1871 10229 1905
rect 10154 1837 10229 1871
rect 10188 1803 10229 1837
rect 10154 1779 10229 1803
rect 9155 1723 9171 1728
rect 9205 1723 9221 1728
rect 10195 1742 10229 1779
rect 9205 1694 9227 1723
rect 9189 1689 9227 1694
rect 9155 1670 9221 1689
rect 10195 1670 10229 1708
rect 8497 1600 8563 1634
rect 8597 1600 8663 1634
rect 8463 1560 8697 1600
rect 10195 1598 10229 1636
rect 12078 2241 12112 2249
rect 12078 2173 12112 2177
rect 12078 2067 12112 2071
rect 12078 1995 12112 2003
rect 12078 1923 12112 1935
rect 12078 1851 12112 1867
rect 12078 1765 12112 1799
rect 12078 1697 12112 1708
rect 12078 1629 12112 1636
rect 8497 1526 8563 1560
rect 8597 1526 8663 1560
rect 8463 1487 8697 1526
rect 8497 1453 8563 1487
rect 8597 1453 8663 1487
rect 8463 1414 8697 1453
rect 8497 1380 8563 1414
rect 8597 1380 8663 1414
rect 8463 1341 8697 1380
rect 8497 1307 8563 1341
rect 8597 1307 8663 1341
rect 8463 1268 8697 1307
rect 8497 1234 8563 1268
rect 8597 1234 8663 1268
rect 8463 1221 8697 1234
rect 12078 1561 12112 1564
rect 12078 1493 12112 1527
rect 12078 1426 12112 1459
rect 12078 1425 12080 1426
rect 12112 1391 12114 1392
rect 12078 1357 12114 1391
rect 12112 1351 12114 1357
rect 12078 1317 12080 1323
rect 12078 1289 12114 1317
rect 12112 1276 12114 1289
rect 12078 1242 12080 1255
rect 12078 1221 12114 1242
rect 12112 1201 12114 1221
rect 12078 1167 12080 1187
rect 12078 1153 12114 1167
rect 12112 1126 12114 1153
rect 12078 1092 12080 1119
rect 12078 1085 12114 1092
rect 12112 1051 12114 1085
rect 12078 1017 12080 1051
rect 17 1002 83 1008
rect -17 968 83 1002
rect 17 934 83 968
rect -17 900 83 934
rect 17 866 83 900
rect -17 832 83 866
rect 17 819 83 832
rect 12112 983 12114 1017
rect 12078 976 12114 983
rect 12078 949 12080 976
rect 12112 915 12114 942
rect 12078 901 12114 915
rect 12078 881 12080 901
rect 12112 847 12114 867
rect 12078 826 12114 847
rect 17 814 661 819
rect 17 810 10605 814
rect 17 798 10472 810
rect -17 781 10472 798
rect -17 747 121 781
rect 155 747 189 781
rect 227 747 257 781
rect 299 747 325 781
rect 371 747 393 781
rect 443 747 461 781
rect 515 747 529 781
rect 587 747 597 781
rect 659 747 665 781
rect 731 747 733 781
rect 767 747 769 781
rect 835 747 841 781
rect 903 747 913 781
rect 971 747 985 781
rect 1039 747 1057 781
rect 1107 747 1129 781
rect 1175 747 1201 781
rect 1243 747 1273 781
rect 1311 747 1345 781
rect 1379 747 1413 781
rect 1451 747 1481 781
rect 1523 747 1549 781
rect 1595 747 1617 781
rect 1667 747 1685 781
rect 1739 747 1753 781
rect 1811 747 1821 781
rect 1883 747 1889 781
rect 1955 747 1957 781
rect 1991 747 1993 781
rect 2059 747 2065 781
rect 2127 747 2137 781
rect 2195 747 2209 781
rect 2263 747 2281 781
rect 2331 747 2353 781
rect 2399 747 2425 781
rect 2467 747 2497 781
rect 2535 747 2569 781
rect 2603 747 2637 781
rect 2675 747 2705 781
rect 2747 747 2773 781
rect 2819 747 2841 781
rect 2891 747 2909 781
rect 2963 747 2977 781
rect 3035 747 3045 781
rect 3107 747 3113 781
rect 3179 747 3181 781
rect 3215 747 3217 781
rect 3283 747 3289 781
rect 3351 747 3361 781
rect 3419 747 3433 781
rect 3487 747 3505 781
rect 3555 747 3577 781
rect 3623 747 3649 781
rect 3691 747 3721 781
rect 3759 747 3793 781
rect 3827 747 3861 781
rect 3899 747 3929 781
rect 3971 747 3997 781
rect 4043 747 4065 781
rect 4115 747 4133 781
rect 4187 747 4201 781
rect 4259 747 4269 781
rect 4331 747 4337 781
rect 4403 747 4405 781
rect 4439 747 4441 781
rect 4507 747 4513 781
rect 4575 747 4585 781
rect 4643 747 4657 781
rect 4711 747 4729 781
rect 4779 747 4801 781
rect 4847 747 4873 781
rect 4915 747 4945 781
rect 4983 747 5017 781
rect 5051 747 5085 781
rect 5123 747 5153 781
rect 5195 747 5221 781
rect 5267 747 5289 781
rect 5339 747 5357 781
rect 5411 747 5425 781
rect 5483 747 5493 781
rect 5555 747 5561 781
rect 5627 747 5629 781
rect 5663 747 5665 781
rect 5731 747 5737 781
rect 5799 747 5809 781
rect 5867 747 5881 781
rect 5935 747 5953 781
rect 6003 747 6025 781
rect 6071 747 6097 781
rect 6139 747 6169 781
rect 6207 747 6241 781
rect 6275 747 6309 781
rect 6347 747 6377 781
rect 6419 747 6445 781
rect 6491 747 6513 781
rect 6563 747 6581 781
rect 6635 747 6649 781
rect 6707 747 6717 781
rect 6779 747 6785 781
rect 6851 747 6853 781
rect 6887 747 6889 781
rect 6955 747 6961 781
rect 7023 747 7033 781
rect 7091 747 7105 781
rect 7159 747 7177 781
rect 7227 747 7249 781
rect 7295 747 7321 781
rect 7363 747 7393 781
rect 7431 747 7465 781
rect 7499 747 7533 781
rect 7571 747 7601 781
rect 7643 747 7669 781
rect 7715 747 7737 781
rect 7787 747 7805 781
rect 7859 747 7873 781
rect 7931 747 7941 781
rect 8003 747 8009 781
rect 8075 747 8077 781
rect 8111 747 8113 781
rect 8179 747 8185 781
rect 8247 747 8257 781
rect 8315 747 8329 781
rect 8383 747 8401 781
rect 8451 747 8473 781
rect 8519 747 8545 781
rect 8587 747 8617 781
rect 8655 747 8689 781
rect 8723 747 8757 781
rect 8795 747 8825 781
rect 8867 747 8893 781
rect 8939 747 8961 781
rect 9011 747 9029 781
rect 9083 747 9097 781
rect 9155 747 9165 781
rect 9227 747 9233 781
rect 9299 747 9301 781
rect 9335 747 9337 781
rect 9403 747 9409 781
rect 9471 747 9481 781
rect 9539 747 9553 781
rect 9607 747 9625 781
rect 9675 747 9697 781
rect 9743 747 9769 781
rect 9811 747 9841 781
rect 9879 747 9913 781
rect 9947 747 9981 781
rect 10019 747 10049 781
rect 10091 747 10117 781
rect 10163 747 10185 781
rect 10235 747 10253 781
rect 10307 747 10321 781
rect 10355 776 10472 781
rect 10506 776 10605 810
rect 12078 813 12080 826
rect 10355 747 10605 776
rect -17 742 10605 747
rect 11671 753 11743 787
rect 11777 753 11824 787
rect 11858 753 11905 787
rect 11939 753 11986 787
rect 12020 779 12078 781
rect 12020 753 12112 779
rect 11671 745 12112 753
rect 11671 742 12078 745
rect -17 714 10519 742
rect 10553 735 10591 742
rect 10505 708 10519 714
rect 10585 708 10591 735
rect 10625 708 10663 742
rect 10697 708 10735 742
rect 10769 708 10807 742
rect 10841 708 10879 742
rect 10913 708 10951 742
rect 10985 708 11023 742
rect 11057 708 11095 742
rect 11129 708 11167 742
rect 11201 708 11239 742
rect 11273 708 11311 742
rect 11345 708 11383 742
rect 11417 708 11455 742
rect 11489 708 11527 742
rect 11561 708 11599 742
rect 11633 711 12078 742
rect 11633 708 12112 711
rect 10505 701 10551 708
rect 10585 701 12112 708
rect 10505 661 12112 701
rect 10505 627 10621 661
rect 10655 627 10692 661
rect 10726 627 10763 661
rect 10797 627 10834 661
rect 10868 627 10905 661
rect 10939 627 10976 661
rect 11010 627 11047 661
rect 11081 627 11118 661
rect 11152 627 11189 661
rect 11223 627 11260 661
rect 11294 627 11331 661
rect 11365 627 11402 661
rect 11436 627 11473 661
rect 11507 627 11544 661
rect 11578 627 11615 661
rect 11649 627 11686 661
rect 11720 627 11757 661
rect 11791 627 11828 661
rect 11862 627 11899 661
rect 11933 627 11970 661
rect 12004 627 12041 661
rect 12075 627 12112 661
rect 10505 623 12112 627
rect 10505 565 12774 623
rect 12104 545 12774 565
rect 12653 487 12774 545
rect 12653 453 12740 487
rect 12653 415 12774 453
rect 12653 381 12740 415
rect 12653 343 12774 381
rect 12653 309 12740 343
rect 12653 -669 12774 309
rect 12494 -708 12774 -669
<< viali >>
rect 333 4437 345 4543
rect 345 4437 787 4543
rect 787 4437 799 4543
rect 12078 4512 12112 4527
rect 12078 4493 12105 4512
rect 12105 4493 12112 4512
rect 12078 4419 12112 4453
rect 12078 4349 12112 4379
rect 12078 4345 12112 4349
rect 8737 4311 8771 4345
rect 8809 4311 8843 4345
rect 12078 4281 12112 4306
rect 12078 4272 12112 4281
rect 12078 4213 12112 4233
rect 12078 4199 12112 4213
rect 12078 4145 12112 4160
rect 12078 4126 12112 4145
rect 7138 3635 7172 3669
rect 7210 3635 7244 3669
rect 7552 3561 7586 3595
rect 7624 3561 7658 3595
rect 7896 3561 7930 3595
rect 7968 3561 8002 3595
rect 8259 3487 8293 3521
rect 8331 3487 8365 3521
rect 8659 3485 8693 3519
rect 8731 3485 8765 3519
rect 9454 3635 9488 3669
rect 9526 3635 9560 3669
rect 9598 3635 9632 3669
rect 9670 3635 9704 3669
rect 9144 3561 9178 3595
rect 9216 3561 9250 3595
rect 9997 3549 10031 3583
rect 10069 3549 10103 3583
rect 10141 3549 10175 3583
rect 9153 3367 9157 3372
rect 9157 3367 9191 3372
rect 9191 3367 9225 3372
rect 9225 3367 9259 3372
rect 9153 3327 9259 3367
rect 9153 3293 9157 3327
rect 9157 3293 9191 3327
rect 9191 3293 9225 3327
rect 9225 3293 9259 3327
rect 9153 3253 9259 3293
rect 9153 3219 9157 3253
rect 9157 3219 9191 3253
rect 9191 3219 9225 3253
rect 9225 3219 9259 3253
rect 9153 3194 9259 3219
rect 11814 3333 11848 3367
rect 11814 3261 11848 3295
rect 11814 3189 11848 3223
rect 12078 3329 12112 3360
rect 12078 3326 12112 3329
rect 12078 3261 12112 3284
rect 12078 3250 12112 3261
rect 12078 3193 12112 3208
rect 12078 3174 12112 3193
rect 12078 3125 12112 3132
rect 12078 3098 12112 3125
rect 12078 3023 12112 3056
rect 12078 3022 12112 3023
rect 12078 2955 12112 2980
rect 12078 2946 12112 2955
rect 12078 2887 12112 2904
rect 12078 2870 12112 2887
rect 12078 2819 12112 2828
rect 12078 2794 12112 2819
rect 12078 2479 12112 2499
rect 12078 2465 12112 2479
rect 12078 2411 12112 2427
rect 12078 2393 12112 2411
rect 12078 2343 12112 2355
rect 12078 2321 12112 2343
rect 12078 2275 12112 2283
rect 3070 2233 3104 2267
rect 3144 2233 3178 2267
rect 3218 2233 3252 2267
rect 3292 2233 3326 2267
rect 3366 2233 3400 2267
rect 3440 2233 3474 2267
rect 3514 2233 3548 2267
rect 3588 2233 3622 2267
rect 3662 2233 3696 2267
rect 3736 2233 3770 2267
rect 3810 2233 3844 2267
rect 3884 2233 3918 2267
rect 3958 2233 3992 2267
rect 4032 2233 4066 2267
rect 4106 2233 4140 2267
rect 4180 2233 4214 2267
rect 4253 2233 4287 2267
rect 4326 2233 4360 2267
rect 4399 2233 4433 2267
rect 4472 2233 4506 2267
rect 4545 2233 4579 2267
rect 4618 2233 4652 2267
rect 9155 1694 9171 1723
rect 9171 1694 9189 1723
rect 9155 1689 9189 1694
rect 9227 1689 9261 1723
rect 10195 1708 10229 1742
rect 10195 1636 10229 1670
rect 10195 1564 10229 1598
rect 12078 2249 12112 2275
rect 12078 2207 12112 2211
rect 12078 2177 12112 2207
rect 12078 2105 12112 2139
rect 12078 2037 12112 2067
rect 12078 2033 12112 2037
rect 12078 1969 12112 1995
rect 12078 1961 12112 1969
rect 12078 1901 12112 1923
rect 12078 1889 12112 1901
rect 12078 1833 12112 1851
rect 12078 1817 12112 1833
rect 12078 1731 12112 1742
rect 12078 1708 12112 1731
rect 12078 1663 12112 1670
rect 12078 1636 12112 1663
rect 12078 1595 12112 1598
rect 12078 1564 12112 1595
rect 12080 1425 12114 1426
rect 12080 1392 12112 1425
rect 12112 1392 12114 1425
rect 12080 1323 12112 1351
rect 12112 1323 12114 1351
rect 12080 1317 12114 1323
rect 12080 1255 12112 1276
rect 12112 1255 12114 1276
rect 12080 1242 12114 1255
rect 8463 1195 8713 1221
rect 8463 1161 8497 1195
rect 8497 1161 8563 1195
rect 8563 1161 8597 1195
rect 8597 1161 8663 1195
rect 8663 1161 8697 1195
rect 8697 1161 8713 1195
rect 8463 1122 8713 1161
rect 8463 1088 8497 1122
rect 8497 1088 8563 1122
rect 8563 1088 8597 1122
rect 8597 1088 8663 1122
rect 8663 1088 8697 1122
rect 8697 1088 8713 1122
rect 8463 1043 8713 1088
rect 12080 1187 12112 1201
rect 12112 1187 12114 1201
rect 12080 1167 12114 1187
rect 12080 1119 12112 1126
rect 12112 1119 12114 1126
rect 12080 1092 12114 1119
rect 12080 1017 12114 1051
rect 12080 949 12114 976
rect 12080 942 12112 949
rect 12112 942 12114 949
rect 12080 881 12114 901
rect 12080 867 12112 881
rect 12112 867 12114 881
rect 121 747 155 781
rect 193 747 223 781
rect 223 747 227 781
rect 265 747 291 781
rect 291 747 299 781
rect 337 747 359 781
rect 359 747 371 781
rect 409 747 427 781
rect 427 747 443 781
rect 481 747 495 781
rect 495 747 515 781
rect 553 747 563 781
rect 563 747 587 781
rect 625 747 631 781
rect 631 747 659 781
rect 697 747 699 781
rect 699 747 731 781
rect 769 747 801 781
rect 801 747 803 781
rect 841 747 869 781
rect 869 747 875 781
rect 913 747 937 781
rect 937 747 947 781
rect 985 747 1005 781
rect 1005 747 1019 781
rect 1057 747 1073 781
rect 1073 747 1091 781
rect 1129 747 1141 781
rect 1141 747 1163 781
rect 1201 747 1209 781
rect 1209 747 1235 781
rect 1273 747 1277 781
rect 1277 747 1307 781
rect 1345 747 1379 781
rect 1417 747 1447 781
rect 1447 747 1451 781
rect 1489 747 1515 781
rect 1515 747 1523 781
rect 1561 747 1583 781
rect 1583 747 1595 781
rect 1633 747 1651 781
rect 1651 747 1667 781
rect 1705 747 1719 781
rect 1719 747 1739 781
rect 1777 747 1787 781
rect 1787 747 1811 781
rect 1849 747 1855 781
rect 1855 747 1883 781
rect 1921 747 1923 781
rect 1923 747 1955 781
rect 1993 747 2025 781
rect 2025 747 2027 781
rect 2065 747 2093 781
rect 2093 747 2099 781
rect 2137 747 2161 781
rect 2161 747 2171 781
rect 2209 747 2229 781
rect 2229 747 2243 781
rect 2281 747 2297 781
rect 2297 747 2315 781
rect 2353 747 2365 781
rect 2365 747 2387 781
rect 2425 747 2433 781
rect 2433 747 2459 781
rect 2497 747 2501 781
rect 2501 747 2531 781
rect 2569 747 2603 781
rect 2641 747 2671 781
rect 2671 747 2675 781
rect 2713 747 2739 781
rect 2739 747 2747 781
rect 2785 747 2807 781
rect 2807 747 2819 781
rect 2857 747 2875 781
rect 2875 747 2891 781
rect 2929 747 2943 781
rect 2943 747 2963 781
rect 3001 747 3011 781
rect 3011 747 3035 781
rect 3073 747 3079 781
rect 3079 747 3107 781
rect 3145 747 3147 781
rect 3147 747 3179 781
rect 3217 747 3249 781
rect 3249 747 3251 781
rect 3289 747 3317 781
rect 3317 747 3323 781
rect 3361 747 3385 781
rect 3385 747 3395 781
rect 3433 747 3453 781
rect 3453 747 3467 781
rect 3505 747 3521 781
rect 3521 747 3539 781
rect 3577 747 3589 781
rect 3589 747 3611 781
rect 3649 747 3657 781
rect 3657 747 3683 781
rect 3721 747 3725 781
rect 3725 747 3755 781
rect 3793 747 3827 781
rect 3865 747 3895 781
rect 3895 747 3899 781
rect 3937 747 3963 781
rect 3963 747 3971 781
rect 4009 747 4031 781
rect 4031 747 4043 781
rect 4081 747 4099 781
rect 4099 747 4115 781
rect 4153 747 4167 781
rect 4167 747 4187 781
rect 4225 747 4235 781
rect 4235 747 4259 781
rect 4297 747 4303 781
rect 4303 747 4331 781
rect 4369 747 4371 781
rect 4371 747 4403 781
rect 4441 747 4473 781
rect 4473 747 4475 781
rect 4513 747 4541 781
rect 4541 747 4547 781
rect 4585 747 4609 781
rect 4609 747 4619 781
rect 4657 747 4677 781
rect 4677 747 4691 781
rect 4729 747 4745 781
rect 4745 747 4763 781
rect 4801 747 4813 781
rect 4813 747 4835 781
rect 4873 747 4881 781
rect 4881 747 4907 781
rect 4945 747 4949 781
rect 4949 747 4979 781
rect 5017 747 5051 781
rect 5089 747 5119 781
rect 5119 747 5123 781
rect 5161 747 5187 781
rect 5187 747 5195 781
rect 5233 747 5255 781
rect 5255 747 5267 781
rect 5305 747 5323 781
rect 5323 747 5339 781
rect 5377 747 5391 781
rect 5391 747 5411 781
rect 5449 747 5459 781
rect 5459 747 5483 781
rect 5521 747 5527 781
rect 5527 747 5555 781
rect 5593 747 5595 781
rect 5595 747 5627 781
rect 5665 747 5697 781
rect 5697 747 5699 781
rect 5737 747 5765 781
rect 5765 747 5771 781
rect 5809 747 5833 781
rect 5833 747 5843 781
rect 5881 747 5901 781
rect 5901 747 5915 781
rect 5953 747 5969 781
rect 5969 747 5987 781
rect 6025 747 6037 781
rect 6037 747 6059 781
rect 6097 747 6105 781
rect 6105 747 6131 781
rect 6169 747 6173 781
rect 6173 747 6203 781
rect 6241 747 6275 781
rect 6313 747 6343 781
rect 6343 747 6347 781
rect 6385 747 6411 781
rect 6411 747 6419 781
rect 6457 747 6479 781
rect 6479 747 6491 781
rect 6529 747 6547 781
rect 6547 747 6563 781
rect 6601 747 6615 781
rect 6615 747 6635 781
rect 6673 747 6683 781
rect 6683 747 6707 781
rect 6745 747 6751 781
rect 6751 747 6779 781
rect 6817 747 6819 781
rect 6819 747 6851 781
rect 6889 747 6921 781
rect 6921 747 6923 781
rect 6961 747 6989 781
rect 6989 747 6995 781
rect 7033 747 7057 781
rect 7057 747 7067 781
rect 7105 747 7125 781
rect 7125 747 7139 781
rect 7177 747 7193 781
rect 7193 747 7211 781
rect 7249 747 7261 781
rect 7261 747 7283 781
rect 7321 747 7329 781
rect 7329 747 7355 781
rect 7393 747 7397 781
rect 7397 747 7427 781
rect 7465 747 7499 781
rect 7537 747 7567 781
rect 7567 747 7571 781
rect 7609 747 7635 781
rect 7635 747 7643 781
rect 7681 747 7703 781
rect 7703 747 7715 781
rect 7753 747 7771 781
rect 7771 747 7787 781
rect 7825 747 7839 781
rect 7839 747 7859 781
rect 7897 747 7907 781
rect 7907 747 7931 781
rect 7969 747 7975 781
rect 7975 747 8003 781
rect 8041 747 8043 781
rect 8043 747 8075 781
rect 8113 747 8145 781
rect 8145 747 8147 781
rect 8185 747 8213 781
rect 8213 747 8219 781
rect 8257 747 8281 781
rect 8281 747 8291 781
rect 8329 747 8349 781
rect 8349 747 8363 781
rect 8401 747 8417 781
rect 8417 747 8435 781
rect 8473 747 8485 781
rect 8485 747 8507 781
rect 8545 747 8553 781
rect 8553 747 8579 781
rect 8617 747 8621 781
rect 8621 747 8651 781
rect 8689 747 8723 781
rect 8761 747 8791 781
rect 8791 747 8795 781
rect 8833 747 8859 781
rect 8859 747 8867 781
rect 8905 747 8927 781
rect 8927 747 8939 781
rect 8977 747 8995 781
rect 8995 747 9011 781
rect 9049 747 9063 781
rect 9063 747 9083 781
rect 9121 747 9131 781
rect 9131 747 9155 781
rect 9193 747 9199 781
rect 9199 747 9227 781
rect 9265 747 9267 781
rect 9267 747 9299 781
rect 9337 747 9369 781
rect 9369 747 9371 781
rect 9409 747 9437 781
rect 9437 747 9443 781
rect 9481 747 9505 781
rect 9505 747 9515 781
rect 9553 747 9573 781
rect 9573 747 9587 781
rect 9625 747 9641 781
rect 9641 747 9659 781
rect 9697 747 9709 781
rect 9709 747 9731 781
rect 9769 747 9777 781
rect 9777 747 9803 781
rect 9841 747 9845 781
rect 9845 747 9875 781
rect 9913 747 9947 781
rect 9985 747 10015 781
rect 10015 747 10019 781
rect 10057 747 10083 781
rect 10083 747 10091 781
rect 10129 747 10151 781
rect 10151 747 10163 781
rect 10201 747 10219 781
rect 10219 747 10235 781
rect 10273 747 10287 781
rect 10287 747 10307 781
rect 12080 813 12114 826
rect 12080 792 12112 813
rect 12112 792 12114 813
rect 11743 753 11777 787
rect 11824 753 11858 787
rect 11905 753 11939 787
rect 11986 753 12020 787
rect 10519 735 10553 742
rect 10519 708 10551 735
rect 10551 708 10553 735
rect 10591 708 10625 742
rect 10663 708 10697 742
rect 10735 708 10769 742
rect 10807 708 10841 742
rect 10879 708 10913 742
rect 10951 708 10985 742
rect 11023 708 11057 742
rect 11095 708 11129 742
rect 11167 708 11201 742
rect 11239 708 11273 742
rect 11311 708 11345 742
rect 11383 708 11417 742
rect 11455 708 11489 742
rect 11527 708 11561 742
rect 11599 708 11633 742
rect 12740 453 12774 487
rect 12740 381 12774 415
rect 12740 309 12774 343
<< metal1 >>
rect -26 4864 35 4867
tri 35 4864 38 4867 sw
rect -26 4818 496 4864
rect -26 4815 51 4818
tri 51 4815 54 4818 nw
rect -26 4563 26 4815
tri 26 4790 51 4815 nw
tri 26 4563 51 4588 sw
rect -26 4543 7986 4563
rect -26 4437 333 4543
rect 799 4437 7986 4543
rect -26 4417 7986 4437
rect 12059 4527 12118 4539
rect 12059 4493 12078 4527
rect 12112 4493 12118 4527
rect 12059 4479 12118 4493
rect 12111 4453 12118 4479
rect 12059 4419 12078 4427
rect 12112 4419 12118 4453
rect -26 3905 26 4417
tri 26 4392 51 4417 nw
rect 12059 4402 12118 4419
rect 12111 4379 12118 4402
rect 8725 4304 8731 4356
rect 8783 4304 8797 4356
rect 8849 4304 8855 4356
rect 12059 4345 12078 4350
rect 12112 4345 12118 4379
rect 12059 4325 12118 4345
rect 12111 4306 12118 4325
rect 12059 4272 12078 4273
rect 12112 4272 12118 4306
rect 12059 4248 12118 4272
tri 10150 4233 10155 4238 se
rect 10155 4233 10207 4238
rect 7138 4232 10207 4233
rect 7138 4205 10155 4232
tri 10130 4199 10136 4205 ne
rect 10136 4199 10155 4205
tri 10136 4194 10141 4199 ne
rect 10141 4194 10155 4199
rect 121 4163 265 4194
tri 10141 4180 10155 4194 ne
rect 7860 4131 7906 4177
rect 9102 4131 9148 4177
rect 10155 4168 10207 4180
rect 10072 4089 10112 4135
rect 10155 4110 10207 4116
rect 12111 4233 12118 4248
rect 12112 4199 12118 4233
rect 12111 4196 12118 4199
rect 12059 4172 12118 4196
rect 12111 4160 12118 4172
rect 12112 4126 12118 4160
rect 12111 4120 12118 4126
rect 12059 4114 12118 4120
rect 7668 4013 7708 4059
rect 5766 3933 5806 3979
rect 5902 3933 5943 3979
tri 26 3905 51 3930 sw
rect -26 3899 12388 3905
rect -26 3847 12059 3899
rect 12111 3847 12388 3899
rect -26 3830 12388 3847
rect -26 3778 12059 3830
rect 12111 3778 12388 3830
rect -26 3761 12388 3778
rect -26 3739 12059 3761
rect -26 3707 1515 3739
tri 1515 3707 1547 3739 nw
tri 1661 3707 1693 3739 ne
rect 1693 3709 12059 3739
rect 12111 3709 12388 3761
rect 1693 3707 12388 3709
rect -26 3703 1511 3707
tri 1511 3703 1515 3707 nw
tri 1693 3703 1697 3707 ne
rect 1697 3703 12388 3707
rect -26 3669 266 3703
tri 266 3669 300 3703 nw
rect -26 3641 238 3669
tri 238 3641 266 3669 nw
rect -26 3635 232 3641
tri 232 3635 238 3641 nw
rect -26 3595 192 3635
tri 192 3595 232 3635 nw
rect 398 3629 435 3675
rect 6875 3669 9716 3675
rect 6927 3635 7138 3669
rect 7172 3635 7210 3669
rect 7244 3635 9454 3669
rect 9488 3635 9526 3669
rect 9560 3635 9598 3669
rect 9632 3635 9670 3669
rect 9704 3635 9716 3669
rect 6927 3629 9086 3635
tri 9086 3629 9092 3635 nw
tri 9285 3629 9291 3635 ne
rect 9291 3629 9716 3635
rect 6875 3605 6927 3617
rect -303 3055 -257 3101
tri -73 2629 -26 2676 se
rect -26 2629 172 3595
tri 172 3575 192 3595 nw
tri 6927 3604 6952 3629 nw
rect 7540 3595 7670 3601
rect 6875 3547 6927 3553
rect 7013 3561 7065 3564
tri 7065 3561 7068 3564 sw
rect 7540 3561 7552 3595
rect 7586 3561 7624 3595
rect 7658 3561 7670 3595
rect 7013 3558 7068 3561
rect 7065 3549 7068 3558
tri 7068 3549 7080 3561 sw
rect 7540 3555 7670 3561
rect 7884 3595 9262 3601
tri 9262 3595 9268 3601 sw
rect 7884 3561 7896 3595
rect 7930 3561 7968 3595
rect 8002 3561 9144 3595
rect 9178 3561 9216 3595
rect 9250 3589 9892 3595
tri 9892 3589 9898 3595 sw
rect 9250 3583 9898 3589
tri 9898 3583 9904 3589 sw
rect 9985 3583 10085 3595
rect 10137 3583 10149 3595
rect 9250 3561 9904 3583
rect 7884 3555 9904 3561
tri 9904 3555 9932 3583 sw
tri 7878 3549 7884 3555 se
rect 7884 3549 8052 3555
tri 8052 3549 8058 3555 nw
tri 9858 3549 9864 3555 ne
rect 9864 3549 9932 3555
tri 9932 3549 9938 3555 sw
rect 9985 3549 9997 3583
rect 10031 3549 10069 3583
rect 10137 3549 10141 3583
rect 7065 3521 7080 3549
tri 7080 3521 7108 3549 sw
tri 7850 3521 7878 3549 se
rect 7878 3521 8024 3549
tri 8024 3521 8052 3549 nw
tri 9864 3527 9886 3549 ne
rect 9886 3527 9938 3549
tri 9938 3527 9960 3549 sw
rect 9985 3543 10085 3549
rect 10137 3543 10149 3549
rect 10201 3543 10207 3595
rect 8247 3521 8377 3527
rect 7065 3520 7108 3521
tri 7108 3520 7109 3521 sw
tri 7849 3520 7850 3521 se
rect 7850 3520 8023 3521
tri 8023 3520 8024 3521 nw
rect 7065 3515 8018 3520
tri 8018 3515 8023 3520 nw
rect 7065 3506 7991 3515
rect 7013 3494 7991 3506
rect 7065 3488 7991 3494
tri 7991 3488 8018 3515 nw
rect 7065 3487 7116 3488
tri 7116 3487 7117 3488 nw
rect 8247 3487 8259 3521
rect 8293 3487 8331 3521
rect 8365 3487 8377 3521
rect 7065 3485 7114 3487
tri 7114 3485 7116 3487 nw
rect 7065 3463 7092 3485
tri 7092 3463 7114 3485 nw
rect 8247 3481 8377 3487
rect 8647 3519 8731 3527
rect 8647 3485 8659 3519
rect 8693 3485 8731 3519
rect 8647 3475 8731 3485
rect 8783 3475 8795 3527
rect 8847 3475 9386 3527
rect 9438 3475 9450 3527
rect 9502 3475 9508 3527
tri 9886 3515 9898 3527 ne
rect 9898 3515 9960 3527
tri 9960 3515 9972 3527 sw
tri 9898 3475 9938 3515 ne
rect 9938 3475 10330 3515
tri 9938 3463 9950 3475 ne
rect 9950 3463 10330 3475
rect 10382 3463 10394 3515
rect 10446 3463 10452 3515
rect 7013 3436 7065 3442
tri 7065 3436 7092 3463 nw
rect 660 3372 10260 3379
rect 660 3194 9153 3372
rect 9259 3367 10260 3372
tri 10260 3367 10272 3379 sw
tri 10504 3367 10516 3379 se
rect 10516 3367 11923 3379
rect 9259 3334 10272 3367
tri 10272 3334 10305 3367 sw
tri 10471 3334 10504 3367 se
rect 10504 3334 11814 3367
rect 9259 3333 11814 3334
rect 11848 3333 11923 3367
rect 9259 3295 11923 3333
rect 9259 3261 11814 3295
rect 11848 3261 11923 3295
rect 9259 3223 11923 3261
rect 9259 3194 11814 3223
rect 660 3189 11814 3194
rect 11848 3189 11923 3223
rect 660 3177 11923 3189
rect 12059 3366 12118 3372
rect 12111 3360 12118 3366
rect 12112 3326 12118 3360
rect 12111 3314 12118 3326
rect 12059 3300 12118 3314
rect 12111 3284 12118 3300
rect 12112 3250 12118 3284
rect 12111 3248 12118 3250
rect 12059 3234 12118 3248
rect 12111 3208 12118 3234
rect 12059 3174 12078 3182
rect 12112 3174 12118 3208
rect 12059 3168 12118 3174
rect 12111 3132 12118 3168
rect 12059 3102 12078 3116
rect 12112 3098 12118 3132
rect 12111 3056 12118 3098
rect 12059 3036 12078 3050
rect 12112 3022 12118 3056
rect 12111 2984 12118 3022
rect 12059 2980 12118 2984
rect 12059 2970 12078 2980
rect 12112 2946 12118 2980
rect 12111 2918 12118 2946
rect 12059 2905 12118 2918
rect 12111 2904 12118 2905
rect 654 2765 12023 2895
rect 12112 2870 12118 2904
rect 12111 2853 12118 2870
rect 12059 2840 12118 2853
rect 12111 2828 12118 2840
rect 12112 2794 12118 2828
rect 12111 2788 12118 2794
rect 12059 2782 12118 2788
rect 11574 2698 11635 2729
rect -136 2588 172 2629
rect -136 2511 95 2588
tri 95 2511 172 2588 nw
rect -136 2499 83 2511
tri 83 2499 95 2511 nw
rect 12059 2505 12118 2511
rect 12111 2499 12118 2505
rect -136 2465 49 2499
tri 49 2465 83 2499 nw
rect 12112 2465 12118 2499
rect -136 2427 11 2465
tri 11 2427 49 2465 nw
rect 12111 2453 12118 2465
rect 12059 2440 12118 2453
rect 12111 2427 12118 2440
rect -136 2426 10 2427
tri 10 2426 11 2427 nw
rect 12112 2393 12118 2427
rect 12111 2388 12118 2393
rect 12059 2375 12118 2388
rect 12111 2355 12118 2375
rect 12059 2321 12078 2323
rect 12112 2321 12118 2355
rect 12059 2311 12118 2321
rect 12111 2283 12118 2311
rect 932 2267 11887 2279
rect 932 2233 3070 2267
rect 3104 2233 3144 2267
rect 3178 2233 3218 2267
rect 3252 2233 3292 2267
rect 3326 2233 3366 2267
rect 3400 2233 3440 2267
rect 3474 2233 3514 2267
rect 3548 2233 3588 2267
rect 3622 2233 3662 2267
rect 3696 2233 3736 2267
rect 3770 2233 3810 2267
rect 3844 2233 3884 2267
rect 3918 2233 3958 2267
rect 3992 2233 4032 2267
rect 4066 2233 4106 2267
rect 4140 2233 4180 2267
rect 4214 2233 4253 2267
rect 4287 2233 4326 2267
rect 4360 2233 4399 2267
rect 4433 2233 4472 2267
rect 4506 2233 4545 2267
rect 4579 2233 4618 2267
rect 4652 2233 11887 2267
rect -459 2165 -257 2207
rect 932 2149 11887 2233
rect 12059 2249 12078 2259
rect 12112 2249 12118 2283
rect 12059 2247 12118 2249
rect 12111 2211 12118 2247
rect 12059 2183 12078 2195
rect 12112 2177 12118 2211
rect 12111 2139 12118 2177
rect 12059 2119 12078 2131
rect 12112 2105 12118 2139
rect 12111 2067 12118 2105
rect 12059 2055 12078 2067
rect 12112 2033 12118 2067
rect 12111 2003 12118 2033
rect 12059 1995 12118 2003
rect 12059 1991 12078 1995
rect 12112 1961 12118 1995
rect 12111 1939 12118 1961
rect 12059 1927 12118 1939
rect 12111 1923 12118 1927
rect 12112 1889 12118 1923
rect 12111 1875 12118 1889
rect 12059 1863 12118 1875
rect 12111 1851 12118 1863
rect 12112 1817 12118 1851
rect 12111 1811 12118 1817
rect 12059 1805 12118 1811
rect 650 1748 12388 1754
rect 650 1742 12059 1748
rect 12111 1742 12388 1748
rect 650 1723 10195 1742
rect 650 1689 9155 1723
rect 9189 1689 9227 1723
rect 9261 1708 10195 1723
rect 10229 1708 12059 1742
rect 12112 1708 12388 1742
rect 9261 1696 12059 1708
rect 12111 1696 12388 1708
rect 9261 1689 12388 1696
rect 650 1679 12388 1689
rect 650 1670 12059 1679
rect 12111 1670 12388 1679
rect -396 1578 -354 1656
rect 650 1636 10195 1670
rect 10229 1636 12059 1670
rect 12112 1636 12388 1670
rect 650 1627 12059 1636
rect 12111 1627 12388 1636
rect 650 1610 12388 1627
rect 650 1598 12059 1610
rect 12111 1598 12388 1610
rect 650 1564 10195 1598
rect 10229 1564 12059 1598
rect 12112 1564 12388 1598
rect 650 1558 12059 1564
rect 12111 1558 12388 1564
rect 650 1552 12388 1558
rect 12059 1432 12120 1438
rect 12111 1426 12120 1432
rect 12114 1392 12120 1426
rect 12111 1380 12120 1392
rect 12059 1366 12120 1380
rect -646 1225 -483 1359
rect 12111 1351 12120 1366
rect 12114 1317 12120 1351
rect 12111 1314 12120 1317
rect 12059 1300 12120 1314
rect 12111 1276 12120 1300
rect 12059 1242 12080 1248
rect 12114 1242 12120 1276
rect 12059 1234 12120 1242
rect 182 1221 8787 1228
rect 182 1043 8463 1221
rect 8713 1043 8787 1221
rect 182 1026 8787 1043
rect 12111 1201 12120 1234
rect 12059 1169 12080 1182
rect 12114 1167 12120 1201
rect 12111 1126 12120 1167
rect 12059 1104 12080 1117
rect 12114 1092 12120 1126
rect 12111 1052 12120 1092
rect 12059 1051 12120 1052
rect 12059 1039 12080 1051
rect 12114 1017 12120 1051
rect 12111 987 12120 1017
rect 12059 976 12120 987
rect 12059 974 12080 976
rect 12114 942 12120 976
rect 12111 922 12120 942
rect 12059 909 12120 922
rect 12111 901 12120 909
tri 12031 867 12059 895 se
rect 12114 867 12120 901
tri 12022 858 12031 867 se
rect 12031 858 12059 867
tri 11594 826 11626 858 se
rect 11626 857 12059 858
rect 12111 857 12120 867
rect 11626 844 12120 857
rect 11626 826 12059 844
rect 12111 826 12120 844
rect 81 781 541 826
rect 81 747 121 781
rect 155 747 193 781
rect 227 747 265 781
rect 299 747 337 781
rect 371 747 409 781
rect 443 747 481 781
rect 515 774 541 781
rect 593 774 606 826
rect 658 781 671 826
rect 723 781 736 826
rect 788 781 801 826
rect 853 781 865 826
rect 917 781 929 826
rect 981 781 993 826
rect 659 774 671 781
rect 731 774 736 781
rect 981 774 985 781
rect 1045 774 1057 826
rect 1109 774 1121 826
rect 1173 774 1185 826
rect 1237 792 12059 826
rect 12114 792 12120 826
rect 1237 787 12120 792
rect 1237 781 11743 787
rect 1237 774 1273 781
rect 515 754 553 774
rect 587 754 625 774
rect 659 754 697 774
rect 731 754 769 774
rect 803 754 841 774
rect 875 754 913 774
rect 947 754 985 774
rect 1019 754 1057 774
rect 1091 754 1129 774
rect 1163 754 1201 774
rect 1235 754 1273 774
rect 515 747 541 754
rect 81 702 541 747
rect 593 702 606 754
rect 659 747 671 754
rect 731 747 736 754
rect 981 747 985 754
rect 658 702 671 747
rect 723 702 736 747
rect 788 702 801 747
rect 853 702 865 747
rect 917 702 929 747
rect 981 702 993 747
rect 1045 702 1057 754
rect 1109 702 1121 754
rect 1173 702 1185 754
rect 1237 747 1273 754
rect 1307 747 1345 781
rect 1379 747 1417 781
rect 1451 747 1489 781
rect 1523 747 1561 781
rect 1595 747 1633 781
rect 1667 747 1705 781
rect 1739 747 1777 781
rect 1811 747 1849 781
rect 1883 747 1921 781
rect 1955 747 1993 781
rect 2027 747 2065 781
rect 2099 747 2137 781
rect 2171 747 2209 781
rect 2243 747 2281 781
rect 2315 747 2353 781
rect 2387 747 2425 781
rect 2459 747 2497 781
rect 2531 747 2569 781
rect 2603 747 2641 781
rect 2675 747 2713 781
rect 2747 747 2785 781
rect 2819 747 2857 781
rect 2891 747 2929 781
rect 2963 747 3001 781
rect 3035 747 3073 781
rect 3107 747 3145 781
rect 3179 747 3217 781
rect 3251 747 3289 781
rect 3323 747 3361 781
rect 3395 747 3433 781
rect 3467 747 3505 781
rect 3539 747 3577 781
rect 3611 747 3649 781
rect 3683 747 3721 781
rect 3755 747 3793 781
rect 3827 747 3865 781
rect 3899 747 3937 781
rect 3971 747 4009 781
rect 4043 747 4081 781
rect 4115 747 4153 781
rect 4187 747 4225 781
rect 4259 747 4297 781
rect 4331 747 4369 781
rect 4403 747 4441 781
rect 4475 747 4513 781
rect 4547 747 4585 781
rect 4619 747 4657 781
rect 4691 747 4729 781
rect 4763 747 4801 781
rect 4835 747 4873 781
rect 4907 747 4945 781
rect 4979 747 5017 781
rect 5051 747 5089 781
rect 5123 747 5161 781
rect 5195 747 5233 781
rect 5267 747 5305 781
rect 5339 747 5377 781
rect 5411 747 5449 781
rect 5483 747 5521 781
rect 5555 747 5593 781
rect 5627 747 5665 781
rect 5699 747 5737 781
rect 5771 747 5809 781
rect 5843 747 5881 781
rect 5915 747 5953 781
rect 5987 747 6025 781
rect 6059 747 6097 781
rect 6131 747 6169 781
rect 6203 747 6241 781
rect 6275 747 6313 781
rect 6347 747 6385 781
rect 6419 747 6457 781
rect 6491 747 6529 781
rect 6563 747 6601 781
rect 6635 747 6673 781
rect 6707 747 6745 781
rect 6779 747 6817 781
rect 6851 747 6889 781
rect 6923 747 6961 781
rect 6995 747 7033 781
rect 7067 747 7105 781
rect 7139 747 7177 781
rect 7211 747 7249 781
rect 7283 747 7321 781
rect 7355 747 7393 781
rect 7427 747 7465 781
rect 7499 747 7537 781
rect 7571 747 7609 781
rect 7643 747 7681 781
rect 7715 747 7753 781
rect 7787 747 7825 781
rect 7859 747 7897 781
rect 7931 747 7969 781
rect 8003 747 8041 781
rect 8075 747 8113 781
rect 8147 747 8185 781
rect 8219 747 8257 781
rect 8291 747 8329 781
rect 8363 747 8401 781
rect 8435 747 8473 781
rect 8507 747 8545 781
rect 8579 747 8617 781
rect 8651 747 8689 781
rect 8723 747 8761 781
rect 8795 747 8833 781
rect 8867 747 8905 781
rect 8939 747 8977 781
rect 9011 747 9049 781
rect 9083 747 9121 781
rect 9155 747 9193 781
rect 9227 747 9265 781
rect 9299 747 9337 781
rect 9371 747 9409 781
rect 9443 747 9481 781
rect 9515 747 9553 781
rect 9587 747 9625 781
rect 9659 747 9697 781
rect 9731 747 9769 781
rect 9803 747 9841 781
rect 9875 747 9913 781
rect 9947 747 9985 781
rect 10019 747 10057 781
rect 10091 747 10129 781
rect 10163 747 10201 781
rect 10235 747 10273 781
rect 10307 753 11743 781
rect 11777 753 11824 787
rect 11858 753 11905 787
rect 11939 753 11986 787
rect 12020 753 12120 787
rect 10307 747 12120 753
rect 1237 742 12120 747
rect 1237 708 10519 742
rect 10553 708 10591 742
rect 10625 708 10663 742
rect 10697 708 10735 742
rect 10769 708 10807 742
rect 10841 708 10879 742
rect 10913 708 10951 742
rect 10985 708 11023 742
rect 11057 708 11095 742
rect 11129 708 11167 742
rect 11201 708 11239 742
rect 11273 708 11311 742
rect 11345 708 11383 742
rect 11417 708 11455 742
rect 11489 708 11527 742
rect 11561 708 11599 742
rect 11633 734 12120 742
rect 11633 708 11711 734
rect 1237 702 11711 708
tri 11711 702 11743 734 nw
rect 12059 493 12111 499
rect 12059 424 12111 441
rect -627 319 -425 361
rect 12059 355 12111 372
rect 12059 297 12111 303
rect 12734 487 12780 499
rect 12734 453 12740 487
rect 12774 453 12780 487
rect 12734 415 12780 453
rect 12734 381 12740 415
rect 12774 381 12780 415
rect 12734 343 12780 381
rect 12734 309 12740 343
rect 12774 309 12780 343
rect 12734 297 12780 309
tri 12304 -720 12310 -714 ne
rect 12310 -720 12316 -668
rect 12368 -720 12380 -668
rect 12432 -720 12438 -668
tri 12438 -720 12444 -714 nw
<< via1 >>
rect 12059 4453 12111 4479
rect 12059 4427 12078 4453
rect 12078 4427 12111 4453
rect 12059 4379 12111 4402
rect 8731 4345 8783 4356
rect 8731 4311 8737 4345
rect 8737 4311 8771 4345
rect 8771 4311 8783 4345
rect 8731 4304 8783 4311
rect 8797 4345 8849 4356
rect 8797 4311 8809 4345
rect 8809 4311 8843 4345
rect 8843 4311 8849 4345
rect 8797 4304 8849 4311
rect 12059 4350 12078 4379
rect 12078 4350 12111 4379
rect 12059 4306 12111 4325
rect 12059 4273 12078 4306
rect 12078 4273 12111 4306
rect 10155 4180 10207 4232
rect 10155 4116 10207 4168
rect 12059 4233 12111 4248
rect 12059 4199 12078 4233
rect 12078 4199 12111 4233
rect 12059 4196 12111 4199
rect 12059 4160 12111 4172
rect 12059 4126 12078 4160
rect 12078 4126 12111 4160
rect 12059 4120 12111 4126
rect 12059 3847 12111 3899
rect 12059 3778 12111 3830
rect 12059 3709 12111 3761
rect 6875 3617 6927 3669
rect 6875 3553 6927 3605
rect 7013 3506 7065 3558
rect 10085 3583 10137 3595
rect 10149 3583 10201 3595
rect 10085 3549 10103 3583
rect 10103 3549 10137 3583
rect 10149 3549 10175 3583
rect 10175 3549 10201 3583
rect 10085 3543 10137 3549
rect 10149 3543 10201 3549
rect 7013 3442 7065 3494
rect 8731 3519 8783 3527
rect 8731 3485 8765 3519
rect 8765 3485 8783 3519
rect 8731 3475 8783 3485
rect 8795 3475 8847 3527
rect 9386 3475 9438 3527
rect 9450 3475 9502 3527
rect 10330 3463 10382 3515
rect 10394 3463 10446 3515
rect 12059 3360 12111 3366
rect 12059 3326 12078 3360
rect 12078 3326 12111 3360
rect 12059 3314 12111 3326
rect 12059 3284 12111 3300
rect 12059 3250 12078 3284
rect 12078 3250 12111 3284
rect 12059 3248 12111 3250
rect 12059 3208 12111 3234
rect 12059 3182 12078 3208
rect 12078 3182 12111 3208
rect 12059 3132 12111 3168
rect 12059 3116 12078 3132
rect 12078 3116 12111 3132
rect 12059 3098 12078 3102
rect 12078 3098 12111 3102
rect 12059 3056 12111 3098
rect 12059 3050 12078 3056
rect 12078 3050 12111 3056
rect 12059 3022 12078 3036
rect 12078 3022 12111 3036
rect 12059 2984 12111 3022
rect 12059 2946 12078 2970
rect 12078 2946 12111 2970
rect 12059 2918 12111 2946
rect 12059 2904 12111 2905
rect 12059 2870 12078 2904
rect 12078 2870 12111 2904
rect 12059 2853 12111 2870
rect 12059 2828 12111 2840
rect 12059 2794 12078 2828
rect 12078 2794 12111 2828
rect 12059 2788 12111 2794
rect 12059 2499 12111 2505
rect 12059 2465 12078 2499
rect 12078 2465 12111 2499
rect 12059 2453 12111 2465
rect 12059 2427 12111 2440
rect 12059 2393 12078 2427
rect 12078 2393 12111 2427
rect 12059 2388 12111 2393
rect 12059 2355 12111 2375
rect 12059 2323 12078 2355
rect 12078 2323 12111 2355
rect 12059 2283 12111 2311
rect 12059 2259 12078 2283
rect 12078 2259 12111 2283
rect 12059 2211 12111 2247
rect 12059 2195 12078 2211
rect 12078 2195 12111 2211
rect 12059 2177 12078 2183
rect 12078 2177 12111 2183
rect 12059 2139 12111 2177
rect 12059 2131 12078 2139
rect 12078 2131 12111 2139
rect 12059 2105 12078 2119
rect 12078 2105 12111 2119
rect 12059 2067 12111 2105
rect 12059 2033 12078 2055
rect 12078 2033 12111 2055
rect 12059 2003 12111 2033
rect 12059 1961 12078 1991
rect 12078 1961 12111 1991
rect 12059 1939 12111 1961
rect 12059 1923 12111 1927
rect 12059 1889 12078 1923
rect 12078 1889 12111 1923
rect 12059 1875 12111 1889
rect 12059 1851 12111 1863
rect 12059 1817 12078 1851
rect 12078 1817 12111 1851
rect 12059 1811 12111 1817
rect 12059 1742 12111 1748
rect 12059 1708 12078 1742
rect 12078 1708 12111 1742
rect 12059 1696 12111 1708
rect 12059 1670 12111 1679
rect 12059 1636 12078 1670
rect 12078 1636 12111 1670
rect 12059 1627 12111 1636
rect 12059 1598 12111 1610
rect 12059 1564 12078 1598
rect 12078 1564 12111 1598
rect 12059 1558 12111 1564
rect 12059 1426 12111 1432
rect 12059 1392 12080 1426
rect 12080 1392 12111 1426
rect 12059 1380 12111 1392
rect 12059 1351 12111 1366
rect 12059 1317 12080 1351
rect 12080 1317 12111 1351
rect 12059 1314 12111 1317
rect 12059 1276 12111 1300
rect 12059 1248 12080 1276
rect 12080 1248 12111 1276
rect 12059 1201 12111 1234
rect 12059 1182 12080 1201
rect 12080 1182 12111 1201
rect 12059 1167 12080 1169
rect 12080 1167 12111 1169
rect 12059 1126 12111 1167
rect 12059 1117 12080 1126
rect 12080 1117 12111 1126
rect 12059 1092 12080 1104
rect 12080 1092 12111 1104
rect 12059 1052 12111 1092
rect 12059 1017 12080 1039
rect 12080 1017 12111 1039
rect 12059 987 12111 1017
rect 12059 942 12080 974
rect 12080 942 12111 974
rect 12059 922 12111 942
rect 12059 901 12111 909
rect 12059 867 12080 901
rect 12080 867 12111 901
rect 12059 857 12111 867
rect 12059 826 12111 844
rect 541 781 593 826
rect 541 774 553 781
rect 553 774 587 781
rect 587 774 593 781
rect 606 781 658 826
rect 671 781 723 826
rect 736 781 788 826
rect 801 781 853 826
rect 865 781 917 826
rect 929 781 981 826
rect 993 781 1045 826
rect 606 774 625 781
rect 625 774 658 781
rect 671 774 697 781
rect 697 774 723 781
rect 736 774 769 781
rect 769 774 788 781
rect 801 774 803 781
rect 803 774 841 781
rect 841 774 853 781
rect 865 774 875 781
rect 875 774 913 781
rect 913 774 917 781
rect 929 774 947 781
rect 947 774 981 781
rect 993 774 1019 781
rect 1019 774 1045 781
rect 1057 781 1109 826
rect 1057 774 1091 781
rect 1091 774 1109 781
rect 1121 781 1173 826
rect 1121 774 1129 781
rect 1129 774 1163 781
rect 1163 774 1173 781
rect 1185 781 1237 826
rect 12059 792 12080 826
rect 12080 792 12111 826
rect 1185 774 1201 781
rect 1201 774 1235 781
rect 1235 774 1237 781
rect 541 747 553 754
rect 553 747 587 754
rect 587 747 593 754
rect 541 702 593 747
rect 606 747 625 754
rect 625 747 658 754
rect 671 747 697 754
rect 697 747 723 754
rect 736 747 769 754
rect 769 747 788 754
rect 801 747 803 754
rect 803 747 841 754
rect 841 747 853 754
rect 865 747 875 754
rect 875 747 913 754
rect 913 747 917 754
rect 929 747 947 754
rect 947 747 981 754
rect 993 747 1019 754
rect 1019 747 1045 754
rect 606 702 658 747
rect 671 702 723 747
rect 736 702 788 747
rect 801 702 853 747
rect 865 702 917 747
rect 929 702 981 747
rect 993 702 1045 747
rect 1057 747 1091 754
rect 1091 747 1109 754
rect 1057 702 1109 747
rect 1121 747 1129 754
rect 1129 747 1163 754
rect 1163 747 1173 754
rect 1121 702 1173 747
rect 1185 747 1201 754
rect 1201 747 1235 754
rect 1235 747 1237 754
rect 1185 702 1237 747
rect 12059 441 12111 493
rect 12059 372 12111 424
rect 12059 303 12111 355
rect 12316 -720 12368 -668
rect 12380 -720 12432 -668
<< metal2 >>
rect 12059 4479 12111 4485
rect 12059 4402 12111 4427
rect 8725 4304 8731 4356
rect 8783 4304 8797 4356
rect 8849 4304 8855 4356
rect 12059 4325 12111 4350
tri 8725 4273 8756 4304 ne
rect 8756 4273 8822 4304
tri 8822 4273 8853 4304 nw
tri 8756 4269 8760 4273 ne
rect 6875 3669 6927 3675
rect 6875 3605 6927 3617
rect 6875 3535 6927 3553
rect 7013 3558 7065 3564
tri 8741 3543 8760 3562 se
rect 8760 3543 8812 4273
tri 8812 4263 8822 4273 nw
rect 12059 4248 12111 4273
rect 10155 4232 10207 4238
rect 10155 4168 10207 4180
tri 10130 3595 10155 3620 se
rect 10155 3595 10207 4116
tri 8812 3543 8837 3568 sw
tri 9447 3543 9456 3552 se
rect 10079 3543 10085 3595
rect 10137 3543 10149 3595
rect 10201 3543 10207 3595
rect 12059 4172 12111 4196
rect 12059 3899 12111 4120
rect 12059 3830 12111 3847
rect 12059 3761 12111 3778
rect 7013 3494 7065 3506
tri 8725 3527 8741 3543 se
rect 8741 3527 8837 3543
tri 8837 3527 8853 3543 sw
tri 9431 3527 9447 3543 se
rect 9447 3527 9456 3543
rect 8725 3475 8731 3527
rect 8783 3475 8795 3527
rect 8847 3475 8853 3527
rect 9380 3475 9386 3527
rect 9438 3475 9450 3527
rect 9502 3475 9508 3527
tri 9431 3463 9443 3475 ne
rect 9443 3463 9456 3475
tri 9443 3450 9456 3463 ne
rect 10324 3463 10330 3515
rect 10382 3463 10394 3515
rect 10446 3463 10452 3515
tri 10324 3450 10337 3463 ne
rect 10337 3450 10405 3463
rect 7013 3436 7065 3442
tri 10337 3438 10349 3450 ne
rect 10349 3438 10405 3450
tri 10405 3438 10430 3463 nw
tri 10315 3055 10349 3089 se
rect 10349 3055 10400 3438
tri 10400 3433 10405 3438 nw
rect 12059 3366 12111 3709
rect 12059 3300 12111 3314
rect 12059 3234 12111 3248
rect 12059 3168 12111 3182
rect 11114 3090 11161 3142
rect 12059 3102 12111 3116
rect 12059 3036 12111 3050
rect 12059 2970 12111 2984
rect 12059 2905 12111 2918
rect 12059 2840 12111 2853
rect 10622 2685 10680 2734
rect 12059 2505 12111 2788
rect 12059 2440 12111 2453
rect 12059 2375 12111 2388
rect 12059 2311 12111 2323
rect 12059 2247 12111 2259
rect 12059 2183 12111 2195
rect 11951 2020 11994 2171
rect 12059 2119 12111 2131
rect 12059 2055 12111 2067
rect 12059 1991 12111 2003
rect 12059 1927 12111 1939
rect 12059 1863 12111 1875
rect 12059 1748 12111 1811
rect 12059 1679 12111 1696
rect 12059 1610 12111 1627
rect 12059 1432 12111 1558
rect 12059 1366 12111 1380
rect 12059 1300 12111 1314
rect 12059 1234 12111 1248
rect 12059 1169 12111 1182
rect 12059 1104 12111 1117
rect 12059 1039 12111 1052
rect 12059 974 12111 987
rect 12059 909 12111 922
rect 12059 844 12111 857
rect 535 774 541 826
rect 593 774 606 826
rect 658 774 671 826
rect 723 774 736 826
rect 788 774 801 826
rect 853 774 865 826
rect 917 774 929 826
rect 981 774 993 826
rect 1045 774 1057 826
rect 1109 774 1121 826
rect 1173 774 1185 826
rect 1237 774 1243 826
rect 535 754 1243 774
rect 535 702 541 754
rect 593 702 606 754
rect 658 702 671 754
rect 723 702 736 754
rect 788 702 801 754
rect 853 702 865 754
rect 917 702 929 754
rect 981 702 993 754
rect 1045 702 1057 754
rect 1109 702 1121 754
rect 1173 702 1185 754
rect 1237 702 1243 754
rect 12059 493 12111 792
rect 12059 424 12111 441
rect 12059 355 12111 372
rect 12059 -92 12111 303
tri 12111 -92 12114 -89 sw
rect 12059 -111 12114 -92
tri 12059 -166 12114 -111 ne
tri 12114 -166 12188 -92 sw
tri 12114 -240 12188 -166 ne
tri 12188 -240 12262 -166 sw
tri 12188 -314 12262 -240 ne
tri 12262 -314 12336 -240 sw
tri 12262 -388 12336 -314 ne
tri 12336 -388 12410 -314 sw
tri 12336 -410 12358 -388 ne
tri 12330 -668 12358 -640 se
rect 12358 -668 12410 -388
tri 12410 -668 12438 -640 sw
rect 12310 -720 12316 -668
rect 12368 -720 12380 -668
rect 12432 -720 12438 -668
use sky130_fd_io__com_pdpredrvr_strong_slowv2  sky130_fd_io__com_pdpredrvr_strong_slowv2_0
timestamp 1663361622
transform -1 0 9387 0 1 2797
box 0 0 872 1568
use sky130_fd_io__com_pdpredrvr_weakv2  sky130_fd_io__com_pdpredrvr_weakv2_0
timestamp 1663361622
transform -1 0 8515 0 1 2797
box -85 8 809 1568
use sky130_fd_io__com_pupredrvr_strong_slowv2  sky130_fd_io__com_pupredrvr_strong_slowv2_0
timestamp 1663361622
transform -1 0 10215 0 1 2797
box -93 0 949 1605
use sky130_fd_io__feas_com_pupredrvr_weak  sky130_fd_io__feas_com_pupredrvr_weak_0
timestamp 1663361622
transform -1 0 7791 0 1 2798
box 21 7 731 1967
use sky130_fd_io__gpio_pupredrvr_strongv2  sky130_fd_io__gpio_pupredrvr_strongv2_0
timestamp 1663361622
transform 1 0 66 0 1 2133
box -66 7 7278 2632
use sky130_fd_io__gpiov2_pdpredrvr_strong  sky130_fd_io__gpiov2_pdpredrvr_strong_0
timestamp 1663361622
transform 1 0 660 0 1 906
box -1618 -706 11544 3924
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1663361622
transform 1 0 7138 0 1 3635
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1663361622
transform -1 0 9250 0 1 3561
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1663361622
transform -1 0 8002 0 1 3561
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1663361622
transform 1 0 8659 0 1 3485
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1663361622
transform -1 0 10175 0 1 3549
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1663361622
transform 0 -1 12112 1 0 1564
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1663361622
transform 0 1 10195 -1 0 1742
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1663361622
transform 1 0 9454 0 1 3635
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_0
timestamp 1663361622
transform 1 0 9153 0 -1 3372
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808266  sky130_fd_pr__via_l1m1__example_55959141808266_0
timestamp 1663361622
transform -1 0 8713 0 -1 1221
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808267  sky130_fd_pr__via_l1m1__example_55959141808267_0
timestamp 1663361622
transform 0 -1 799 -1 0 4543
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1663361622
transform 0 1 6875 1 0 3547
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1663361622
transform 0 -1 10207 -1 0 4238
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1663361622
transform 1 0 10079 0 -1 3595
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1663361622
transform -1 0 9508 0 -1 3527
box 0 0 1 1
<< labels >>
flabel metal2 s 11114 3090 11161 3142 3 FreeSans 300 0 0 0 PD_H[3]
port 1 nsew
flabel metal2 s 10622 2685 10680 2734 3 FreeSans 300 0 0 0 PD_H[2]
port 2 nsew
flabel metal2 s 11951 2020 11994 2171 3 FreeSans 520 180 0 0 PDEN_H_N[1]
port 3 nsew
flabel metal2 s 6875 3535 6927 3587 3 FreeSans 300 0 0 0 DRVHI_H
port 4 nsew
flabel metal2 s 10360 3463 10407 3515 7 FreeSans 300 180 0 0 DRVLO_H_N
port 5 nsew
flabel metal1 s -646 1225 -483 1359 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 5902 3933 5943 3979 3 FreeSans 300 0 0 0 PU_H_N[3]
port 7 nsew
flabel metal1 s 5766 3933 5806 3979 7 FreeSans 300 0 0 0 PU_H_N[2]
port 8 nsew
flabel metal1 s 10072 4089 10112 4135 3 FreeSans 300 0 0 0 PU_H_N[1]
port 9 nsew
flabel metal1 s 7668 4013 7708 4059 3 FreeSans 300 0 0 0 PU_H_N[0]
port 10 nsew
flabel metal1 s 9102 4131 9148 4177 3 FreeSans 300 0 0 0 PD_H[1]
port 11 nsew
flabel metal1 s 7860 4131 7906 4177 3 FreeSans 300 0 0 0 PD_H[0]
port 12 nsew
flabel metal1 s 11574 2698 11635 2729 3 FreeSans 520 0 0 0 PD_H[4]
port 13 nsew
flabel metal1 s -303 3055 -257 3101 3 FreeSans 300 0 0 0 SLOW_H
port 14 nsew
flabel metal1 s 121 4163 265 4194 3 FreeSans 520 0 0 0 PUEN_H[1]
port 15 nsew
flabel metal1 s 7550 3563 7644 3594 3 FreeSans 520 0 0 0 PUEN_H[0]
port 16 nsew
flabel metal1 s 8278 3492 8364 3516 3 FreeSans 520 0 0 0 PDEN_H_N[0]
port 17 nsew
flabel metal1 s 11881 3177 11923 3379 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 12346 3703 12388 3905 7 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 7926 4417 7963 4563 7 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 11972 2765 12014 2895 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 11845 2149 11887 2279 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 8745 1026 8787 1228 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 12346 1552 12388 1754 7 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 666 1552 708 1754 3 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 182 1026 224 1228 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 932 2149 974 2279 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 654 2765 696 2895 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 0 4417 37 4563 3 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 0 3703 42 3905 3 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 681 3177 723 3379 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 398 3629 435 3675 7 FreeSans 300 180 0 0 SLOW_H_N
port 20 nsew
flabel metal1 s -396 1578 -354 1656 3 FreeSans 520 90 0 0 I2C_MODE_H_N
port 21 nsew
flabel metal1 s -627 319 -425 361 3 FreeSans 300 90 0 0 VCC_IO
port 19 nsew
flabel metal1 s -459 2165 -257 2207 3 FreeSans 300 90 0 0 VCC_IO
port 19 nsew
flabel comment s 10763 879 10763 879 0 FreeSans 440 0 0 0 LIJUMPER_OK
flabel comment s 560 2408 560 2408 0 FreeSans 300 0 0 0 CONDIODE
flabel comment s 10707 3958 10707 3958 0 FreeSans 300 0 0 0 PDEN_H_N1
flabel comment s 9376 4044 9376 4044 0 FreeSans 300 0 0 0 PDEN_H_N1
flabel comment s 7497 3968 7497 3968 0 FreeSans 300 0 0 0 PDEN_H_N1
flabel comment s 7988 3576 7988 3576 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 9129 3579 9129 3579 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 10392 3490 10392 3490 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 8484 4228 8484 4228 0 FreeSans 300 0 0 0 PUEN_H1
flabel comment s 9328 4228 9328 4228 0 FreeSans 300 0 0 0 PUEN_H1
<< properties >>
string GDS_END 49138340
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 49061462
<< end >>
