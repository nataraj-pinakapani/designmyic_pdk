magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 11 11 11 11 6 C0
port 1 nsew
rlabel  s 11 10 11 11 6 C0
port 1 nsew
rlabel  s 11 10 11 10 6 C0
port 1 nsew
rlabel  s 11 9 11 10 6 C0
port 1 nsew
rlabel  s 11 9 11 9 6 C0
port 1 nsew
rlabel  s 11 8 11 9 6 C0
port 1 nsew
rlabel  s 11 8 11 8 6 C0
port 1 nsew
rlabel  s 11 7 11 7 6 C0
port 1 nsew
rlabel  s 11 6 11 7 6 C0
port 1 nsew
rlabel  s 11 6 11 6 6 C0
port 1 nsew
rlabel  s 11 6 11 6 6 C0
port 1 nsew
rlabel  s 11 5 11 5 6 C0
port 1 nsew
rlabel  s 11 4 11 5 6 C0
port 1 nsew
rlabel  s 11 4 11 4 6 C0
port 1 nsew
rlabel  s 11 3 11 4 6 C0
port 1 nsew
rlabel  s 11 3 11 3 6 C0
port 1 nsew
rlabel  s 11 2 11 2 6 C0
port 1 nsew
rlabel  s 11 1 11 2 6 C0
port 1 nsew
rlabel  s 11 1 11 1 6 C0
port 1 nsew
rlabel  s 11 0 11 1 8 C0
port 1 nsew
rlabel  s 6 11 11 11 6 C0
port 1 nsew
rlabel  s 6 10 11 10 6 C0
port 1 nsew
rlabel  s 6 10 11 10 6 C0
port 1 nsew
rlabel  s 6 9 11 9 6 C0
port 1 nsew
rlabel  s 6 9 11 9 6 C0
port 1 nsew
rlabel  s 6 8 11 8 6 C0
port 1 nsew
rlabel  s 6 7 11 8 6 C0
port 1 nsew
rlabel  s 6 7 11 7 6 C0
port 1 nsew
rlabel  s 6 6 11 6 6 C0
port 1 nsew
rlabel  s 6 5 11 6 6 C0
port 1 nsew
rlabel  s 6 5 11 5 6 C0
port 1 nsew
rlabel  s 6 4 11 4 6 C0
port 1 nsew
rlabel  s 6 4 11 4 6 C0
port 1 nsew
rlabel  s 6 3 11 3 6 C0
port 1 nsew
rlabel  s 6 2 11 3 6 C0
port 1 nsew
rlabel  s 6 2 11 2 6 C0
port 1 nsew
rlabel  s 6 1 11 1 6 C0
port 1 nsew
rlabel  s 6 1 11 1 6 C0
port 1 nsew
rlabel  s 6 11 11 12 6 C0
port 1 nsew
rlabel  s 6 0 11 0 8 C0
port 1 nsew
rlabel  s 0 11 5 12 6 C0
port 1 nsew
rlabel  s 0 11 0 11 4 C0
port 1 nsew
rlabel  s 0 11 5 11 6 C0
port 1 nsew
rlabel  s 0 10 0 11 4 C0
port 1 nsew
rlabel  s 0 10 5 10 6 C0
port 1 nsew
rlabel  s 0 10 0 10 4 C0
port 1 nsew
rlabel  s 0 10 5 10 6 C0
port 1 nsew
rlabel  s 0 9 0 10 4 C0
port 1 nsew
rlabel  s 0 9 5 9 6 C0
port 1 nsew
rlabel  s 0 9 0 9 4 C0
port 1 nsew
rlabel  s 0 9 5 9 6 C0
port 1 nsew
rlabel  s 0 8 0 9 4 C0
port 1 nsew
rlabel  s 0 8 5 8 6 C0
port 1 nsew
rlabel  s 0 8 0 8 4 C0
port 1 nsew
rlabel  s 0 7 5 8 6 C0
port 1 nsew
rlabel  s 0 7 0 7 4 C0
port 1 nsew
rlabel  s 0 7 5 7 6 C0
port 1 nsew
rlabel  s 0 6 0 7 4 C0
port 1 nsew
rlabel  s 0 6 5 6 6 C0
port 1 nsew
rlabel  s 0 6 0 6 4 C0
port 1 nsew
rlabel  s 0 6 0 6 4 C0
port 1 nsew
rlabel  s 0 5 5 6 6 C0
port 1 nsew
rlabel  s 0 5 0 5 4 C0
port 1 nsew
rlabel  s 0 5 5 5 6 C0
port 1 nsew
rlabel  s 0 4 0 5 4 C0
port 1 nsew
rlabel  s 0 4 5 4 6 C0
port 1 nsew
rlabel  s 0 4 0 4 4 C0
port 1 nsew
rlabel  s 0 4 5 4 6 C0
port 1 nsew
rlabel  s 0 3 0 4 4 C0
port 1 nsew
rlabel  s 0 3 5 3 6 C0
port 1 nsew
rlabel  s 0 3 0 3 4 C0
port 1 nsew
rlabel  s 0 2 5 3 6 C0
port 1 nsew
rlabel  s 0 2 0 2 4 C0
port 1 nsew
rlabel  s 0 2 5 2 6 C0
port 1 nsew
rlabel  s 0 1 0 2 4 C0
port 1 nsew
rlabel  s 0 1 5 1 6 C0
port 1 nsew
rlabel  s 0 1 0 1 4 C0
port 1 nsew
rlabel  s 0 1 5 1 6 C0
port 1 nsew
rlabel  s 0 0 0 1 2 C0
port 1 nsew
rlabel  s 0 0 5 0 8 C0
port 1 nsew
rlabel  s 6 11 6 12 6 C1
port 2 nsew
rlabel  s 6 0 6 0 8 C1
port 2 nsew
rlabel  s 6 11 6 11 6 C1
port 2 nsew
rlabel  s 6 10 6 11 6 C1
port 2 nsew
rlabel  s 6 10 6 10 6 C1
port 2 nsew
rlabel  s 6 9 6 9 6 C1
port 2 nsew
rlabel  s 6 8 6 9 6 C1
port 2 nsew
rlabel  s 6 8 6 8 6 C1
port 2 nsew
rlabel  s 6 7 6 8 6 C1
port 2 nsew
rlabel  s 6 7 6 7 6 C1
port 2 nsew
rlabel  s 6 6 6 7 6 C1
port 2 nsew
rlabel  s 6 5 6 6 6 C1
port 2 nsew
rlabel  s 6 5 6 5 6 C1
port 2 nsew
rlabel  s 6 4 6 4 6 C1
port 2 nsew
rlabel  s 6 3 6 4 6 C1
port 2 nsew
rlabel  s 6 3 6 3 6 C1
port 2 nsew
rlabel  s 6 2 6 3 6 C1
port 2 nsew
rlabel  s 6 2 6 2 6 C1
port 2 nsew
rlabel  s 6 1 6 2 6 C1
port 2 nsew
rlabel  s 6 1 6 1 6 C1
port 2 nsew
rlabel  s 0 11 11 11 6 C1
port 2 nsew
rlabel  s 0 11 11 11 6 C1
port 2 nsew
rlabel  s 0 10 11 10 6 C1
port 2 nsew
rlabel  s 0 9 11 10 6 C1
port 2 nsew
rlabel  s 0 9 11 9 6 C1
port 2 nsew
rlabel  s 0 8 11 8 6 C1
port 2 nsew
rlabel  s 0 8 11 8 6 C1
port 2 nsew
rlabel  s 0 7 11 7 6 C1
port 2 nsew
rlabel  s 0 7 11 7 6 C1
port 2 nsew
rlabel  s 0 5 11 5 6 C1
port 2 nsew
rlabel  s 0 4 11 5 6 C1
port 2 nsew
rlabel  s 0 4 11 4 6 C1
port 2 nsew
rlabel  s 0 3 11 3 6 C1
port 2 nsew
rlabel  s 0 3 11 3 6 C1
port 2 nsew
rlabel  s 0 2 11 2 6 C1
port 2 nsew
rlabel  s 0 2 11 2 6 C1
port 2 nsew
rlabel  s 0 1 11 1 6 C1
port 2 nsew
rlabel  s 0 0 11 1 8 C1
port 2 nsew
rlabel  s 0 6 11 6 6 C1
port 2 nsew
rlabel  s 0 6 11 6 6 C1
port 2 nsew
rlabel  s 0 6 11 6 6 C1
port 2 nsew
rlabel metal_blue s 6 6 6 7 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 11 12
string LEFview TRUE
string gencell sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield
string library sky130
string parameter m=1
<< end >>
