magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 53 75 56 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 48 75 51 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 9 1 14 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 9 75 14 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 9 1 13 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 9 75 13 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 69 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 64 1 68 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 68 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel 
 s 0 52 24 53 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 1 48 24 48 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 1 56 24 57 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 1 37 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 50 37 74 40 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 50 48 74 48 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 50 52 74 53 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 50 56 74 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 37 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 24 48 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 52 24 53 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 56 24 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 50 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 50 48 75 48 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 50 52 75 53 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 50 56 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 1 57 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 48 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 56 74 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 53 74 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 52 74 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 52 74 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 48 74 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 40 74 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 39 74 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 39 74 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 39 74 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 38 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 38 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 53 74 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 52 74 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 52 74 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 40 74 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 39 74 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 39 74 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 39 74 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 38 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 38 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 56 74 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 48 74 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 53 73 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 52 73 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 52 73 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 40 73 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 39 73 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 39 73 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 39 73 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 56 73 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 48 73 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 53 73 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 52 73 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 52 73 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 40 73 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 39 73 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 39 73 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 39 73 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 56 73 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 48 73 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 53 73 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 52 73 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 52 73 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 40 73 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 73 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 73 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 73 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 56 73 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 48 73 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 53 72 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 52 72 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 52 72 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 40 72 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 72 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 72 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 72 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 56 72 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 48 72 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 53 72 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 52 72 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 52 72 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 40 72 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 72 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 72 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 39 72 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 56 72 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 48 72 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 53 71 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 52 71 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 52 71 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 40 71 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 39 71 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 39 71 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 39 71 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 56 71 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 48 71 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 53 71 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 52 71 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 52 71 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 40 71 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 39 71 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 39 71 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 39 71 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 56 71 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 48 71 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 53 71 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 52 71 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 52 71 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 40 71 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 71 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 71 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 71 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 56 71 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 48 71 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 53 70 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 52 70 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 52 70 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 40 70 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 70 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 70 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 70 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 56 70 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 48 70 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 53 70 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 52 70 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 52 70 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 40 70 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 70 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 70 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 39 70 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 56 70 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 48 70 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 53 69 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 52 69 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 52 69 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 40 69 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 39 69 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 39 69 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 39 69 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 56 69 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 48 69 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 53 69 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 52 69 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 52 69 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 40 69 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 39 69 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 39 69 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 39 69 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 56 69 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 48 69 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 53 69 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 52 69 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 52 69 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 40 69 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 69 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 69 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 69 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 56 69 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 48 69 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 53 68 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 52 68 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 52 68 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 40 68 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 68 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 68 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 68 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 56 68 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 48 68 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 53 68 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 52 68 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 52 68 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 40 68 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 68 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 68 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 39 68 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 56 68 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 48 68 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 53 67 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 52 67 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 52 67 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 40 67 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 39 67 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 39 67 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 39 67 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 56 67 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 48 67 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 53 67 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 52 67 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 52 67 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 40 67 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 39 67 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 39 67 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 39 67 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 56 67 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 48 67 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 53 67 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 52 67 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 52 67 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 40 67 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 39 67 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 39 67 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 39 67 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 56 66 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 48 66 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 53 66 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 52 66 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 52 66 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 40 66 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 39 66 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 39 66 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 39 66 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 38 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 38 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 56 66 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 48 66 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 53 66 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 52 66 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 52 66 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 40 66 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 66 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 66 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 66 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 56 66 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 48 66 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 53 65 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 52 65 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 52 65 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 40 65 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 65 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 65 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 65 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 56 65 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 48 65 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 53 65 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 52 65 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 52 65 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 40 65 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 65 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 65 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 39 65 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 56 65 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 48 65 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 53 64 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 52 64 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 52 64 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 40 64 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 39 64 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 39 64 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 39 64 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 56 64 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 48 64 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 53 64 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 52 64 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 52 64 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 40 64 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 39 64 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 39 64 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 39 64 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 56 64 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 48 64 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 53 64 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 52 64 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 52 64 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 40 64 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 64 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 64 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 64 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 56 64 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 48 64 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 53 63 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 52 63 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 52 63 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 40 63 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 63 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 63 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 63 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 56 63 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 48 63 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 53 63 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 52 63 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 52 63 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 40 63 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 63 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 63 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 39 63 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 56 63 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 48 63 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 53 62 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 52 62 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 52 62 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 40 62 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 39 62 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 39 62 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 39 62 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 56 62 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 48 62 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 53 62 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 52 62 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 52 62 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 40 62 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 39 62 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 39 62 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 39 62 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 56 62 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 48 62 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 53 62 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 52 62 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 52 62 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 40 62 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 62 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 62 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 62 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 56 62 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 48 62 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 53 61 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 52 61 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 52 61 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 40 61 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 61 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 61 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 61 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 56 61 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 48 61 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 53 61 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 52 61 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 52 61 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 40 61 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 61 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 61 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 39 61 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 56 61 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 48 61 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 53 60 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 52 60 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 52 60 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 40 60 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 39 60 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 39 60 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 39 60 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 56 60 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 48 60 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 53 60 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 52 60 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 52 60 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 40 60 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 39 60 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 39 60 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 39 60 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 56 60 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 48 60 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 53 60 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 52 60 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 52 60 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 40 60 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 60 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 60 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 60 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 56 60 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 48 60 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 53 59 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 52 59 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 52 59 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 40 59 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 59 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 59 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 59 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 56 59 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 48 59 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 53 59 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 52 59 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 52 59 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 40 59 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 59 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 59 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 39 59 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 56 59 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 48 59 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 53 58 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 52 58 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 52 58 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 40 58 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 39 58 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 39 58 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 39 58 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 56 58 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 48 58 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 53 58 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 52 58 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 52 58 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 40 58 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 39 58 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 39 58 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 39 58 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 56 58 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 48 58 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 53 58 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 52 58 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 52 58 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 40 58 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 58 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 58 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 58 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 56 58 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 48 58 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 53 57 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 52 57 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 52 57 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 40 57 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 57 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 57 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 57 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 56 57 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 48 57 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 53 57 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 52 57 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 52 57 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 40 57 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 57 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 57 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 39 57 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 56 57 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 48 57 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 53 56 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 52 56 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 52 56 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 40 56 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 39 56 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 39 56 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 39 56 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 56 56 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 48 56 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 53 56 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 52 56 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 52 56 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 40 56 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 39 56 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 39 56 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 39 56 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 56 56 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 48 56 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 53 56 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 52 56 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 52 56 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 40 56 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 56 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 56 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 56 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 56 56 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 48 56 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 53 55 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 52 55 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 52 55 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 40 55 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 55 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 55 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 55 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 56 55 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 48 55 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 53 55 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 52 55 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 52 55 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 40 55 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 55 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 55 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 39 55 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 56 55 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 48 55 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 53 54 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 52 54 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 52 54 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 40 54 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 39 54 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 39 54 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 39 54 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 56 54 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 48 54 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 53 54 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 52 54 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 52 54 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 40 54 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 39 54 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 39 54 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 39 54 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 56 54 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 48 54 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 53 54 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 52 54 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 52 54 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 40 54 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 54 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 54 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 54 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 56 54 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 48 54 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 53 53 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 52 53 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 52 53 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 40 53 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 53 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 53 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 53 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 56 53 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 48 53 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 53 53 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 52 53 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 52 53 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 40 53 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 53 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 53 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 39 53 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 56 53 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 48 53 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 53 52 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 52 52 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 52 52 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 40 52 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 39 52 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 39 52 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 39 52 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 56 52 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 48 52 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 53 52 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 52 52 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 52 52 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 40 52 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 39 52 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 39 52 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 39 52 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 56 52 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 48 52 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 53 52 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 52 52 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 52 52 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 40 52 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 39 52 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 39 52 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 39 52 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 56 51 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 48 51 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 53 51 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 52 51 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 52 51 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 40 51 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 39 51 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 39 51 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 39 51 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 38 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 38 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 56 51 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 48 51 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 56 51 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 53 51 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 52 51 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 52 51 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 48 51 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 40 51 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 39 51 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 39 51 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 39 51 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 38 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 38 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 50 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 56 24 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 53 24 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 52 24 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 52 24 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 48 24 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 40 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 39 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 39 24 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 39 24 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 56 24 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 48 24 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 40 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 39 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 39 24 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 39 24 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 53 24 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 52 24 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 52 24 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 40 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 24 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 24 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 24 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 56 24 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 48 24 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 53 23 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 52 23 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 52 23 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 40 23 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 23 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 23 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 23 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 56 23 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 48 23 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 53 23 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 52 23 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 52 23 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 40 23 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 23 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 23 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 39 23 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 56 23 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 48 23 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 53 23 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 52 23 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 52 23 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 40 22 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 39 22 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 39 22 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 39 22 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 56 22 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 48 22 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 53 22 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 52 22 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 52 22 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 40 22 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 39 22 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 39 22 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 39 22 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 56 22 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 48 22 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 53 22 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 52 22 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 52 22 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 40 22 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 22 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 22 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 22 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 56 21 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 48 21 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 53 21 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 52 21 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 52 21 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 40 21 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 21 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 21 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 21 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 56 21 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 48 21 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 53 21 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 52 21 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 52 21 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 40 21 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 21 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 21 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 39 21 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 56 21 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 48 21 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 53 21 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 52 21 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 52 21 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 40 20 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 39 20 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 39 20 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 39 20 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 38 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 38 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 56 20 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 48 20 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 53 20 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 52 20 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 52 20 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 40 20 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 39 20 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 39 20 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 39 20 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 38 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 38 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 56 20 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 48 20 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 53 20 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 52 20 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 52 20 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 40 19 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 39 19 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 39 19 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 39 19 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 56 19 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 48 19 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 53 19 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 52 19 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 52 19 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 40 19 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 39 19 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 39 19 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 39 19 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 56 19 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 48 19 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 53 19 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 52 19 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 52 19 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 40 19 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 19 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 19 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 19 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 56 19 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 48 19 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 53 19 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 52 19 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 52 19 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 40 18 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 18 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 18 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 18 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 56 18 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 48 18 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 53 18 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 52 18 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 52 18 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 40 18 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 18 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 18 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 39 18 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 56 18 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 48 18 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 53 18 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 52 18 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 52 18 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 40 17 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 39 17 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 39 17 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 39 17 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 56 17 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 48 17 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 53 17 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 52 17 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 52 17 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 40 17 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 39 17 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 39 17 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 39 17 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 56 17 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 48 17 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 53 17 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 52 17 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 52 17 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 40 17 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 17 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 17 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 17 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 56 17 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 48 17 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 53 17 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 52 17 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 52 17 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 40 16 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 16 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 16 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 16 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 56 16 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 48 16 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 53 16 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 52 16 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 52 16 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 40 16 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 16 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 16 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 39 16 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 56 16 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 48 16 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 53 16 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 52 16 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 52 16 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 40 15 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 39 15 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 39 15 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 39 15 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 56 15 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 48 15 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 53 15 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 52 15 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 52 15 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 40 15 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 39 15 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 39 15 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 39 15 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 56 15 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 48 15 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 53 15 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 52 15 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 52 15 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 40 15 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 15 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 15 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 15 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 56 15 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 48 15 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 53 15 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 52 15 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 52 15 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 40 14 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 14 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 14 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 14 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 56 14 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 48 14 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 53 14 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 52 14 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 52 14 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 40 14 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 14 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 14 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 39 14 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 56 14 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 48 14 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 53 14 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 52 14 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 52 14 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 40 13 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 39 13 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 39 13 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 39 13 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 56 13 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 48 13 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 53 13 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 52 13 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 52 13 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 40 13 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 39 13 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 39 13 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 39 13 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 56 13 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 48 13 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 53 13 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 52 13 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 52 13 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 40 13 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 13 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 13 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 13 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 56 13 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 48 13 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 53 13 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 52 13 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 52 13 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 40 12 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 12 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 12 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 12 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 56 12 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 48 12 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 53 12 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 52 12 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 52 12 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 40 12 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 12 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 12 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 39 12 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 56 12 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 48 12 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 53 12 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 52 12 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 52 12 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 40 11 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 39 11 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 39 11 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 39 11 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 56 11 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 48 11 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 53 11 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 52 11 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 52 11 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 40 11 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 39 11 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 39 11 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 39 11 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 56 11 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 48 11 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 53 11 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 52 11 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 52 11 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 40 11 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 11 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 11 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 11 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 56 11 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 48 11 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 53 11 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 52 11 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 52 11 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 40 10 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 10 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 10 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 10 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 56 10 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 48 10 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 53 10 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 52 10 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 52 10 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 40 10 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 10 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 10 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 39 10 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 56 10 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 48 10 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 53 10 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 52 10 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 52 10 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 40 9 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 39 9 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 39 9 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 39 9 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 56 9 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 48 9 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 53 9 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 52 9 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 52 9 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 40 9 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 39 9 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 39 9 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 39 9 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 56 9 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 48 9 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 53 9 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 52 9 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 52 9 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 40 9 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 9 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 9 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 9 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 56 9 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 48 9 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 53 9 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 52 9 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 52 9 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 40 8 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 8 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 8 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 8 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 56 8 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 48 8 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 53 8 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 52 8 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 52 8 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 40 8 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 8 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 8 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 39 8 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 56 8 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 48 8 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 53 8 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 52 8 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 52 8 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 40 7 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 39 7 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 39 7 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 39 7 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 56 7 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 48 7 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 53 7 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 52 7 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 52 7 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 40 7 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 39 7 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 39 7 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 39 7 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 56 7 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 48 7 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 53 7 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 52 7 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 52 7 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 40 7 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 7 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 7 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 7 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 56 6 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 48 6 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 53 6 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 52 6 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 52 6 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 40 6 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 6 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 6 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 6 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 56 6 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 48 6 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 53 6 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 52 6 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 52 6 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 40 6 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 6 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 6 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 39 6 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 56 6 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 48 6 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 53 6 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 52 6 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 52 6 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 40 5 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 39 5 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 39 5 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 39 5 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 56 5 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 48 5 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 53 5 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 52 5 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 52 5 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 40 5 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 39 5 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 39 5 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 39 5 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 56 5 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 48 5 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 53 5 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 52 5 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 52 5 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 40 5 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 39 5 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 39 5 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 39 5 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 56 4 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 48 4 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 53 4 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 52 4 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 52 4 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 40 4 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 39 4 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 39 4 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 39 4 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 38 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 38 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 56 4 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 48 4 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 53 4 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 52 4 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 52 4 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 40 4 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 4 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 4 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 4 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 56 4 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 48 4 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 53 4 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 52 4 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 52 4 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 40 3 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 3 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 3 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 3 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 56 3 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 48 3 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 53 3 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 52 3 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 52 3 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 40 3 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 3 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 3 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 39 3 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 56 3 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 48 3 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 53 3 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 52 3 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 52 3 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 40 2 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 39 2 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 39 2 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 39 2 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 56 2 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 48 2 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 53 2 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 52 2 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 52 2 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 40 2 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 39 2 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 39 2 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 39 2 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 56 2 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 48 2 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 53 2 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 52 2 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 52 2 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 40 2 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 39 2 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 39 2 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 39 2 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 56 2 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 48 2 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 53 2 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 52 2 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 52 2 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 40 1 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 39 1 40 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 39 1 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 39 1 39 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 38 1 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 38 1 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 56 1 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 48 1 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 53 1 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 52 1 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 52 1 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 56 1 57 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 48 1 48 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 53 1 53 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 52 1 52 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 52 1 52 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
