magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 11 10 11 11 6 C0
port 1 nsew
rlabel  s 11 9 11 10 6 C0
port 1 nsew
rlabel  s 11 8 11 9 6 C0
port 1 nsew
rlabel  s 11 7 11 8 6 C0
port 1 nsew
rlabel  s 11 5 11 6 6 C0
port 1 nsew
rlabel  s 11 4 11 5 6 C0
port 1 nsew
rlabel  s 11 3 11 4 6 C0
port 1 nsew
rlabel  s 11 2 11 2 6 C0
port 1 nsew
rlabel  s 11 0 11 1 8 C0
port 1 nsew
rlabel  s 6 10 11 10 6 C0
port 1 nsew
rlabel  s 6 9 11 9 6 C0
port 1 nsew
rlabel  s 6 8 11 8 6 C0
port 1 nsew
rlabel  s 6 6 11 7 6 C0
port 1 nsew
rlabel  s 6 5 11 5 6 C0
port 1 nsew
rlabel  s 6 4 11 4 6 C0
port 1 nsew
rlabel  s 6 2 11 3 6 C0
port 1 nsew
rlabel  s 6 1 11 2 6 C0
port 1 nsew
rlabel  s 0 11 11 12 6 C0
port 1 nsew
rlabel  s 0 10 0 11 4 C0
port 1 nsew
rlabel  s 0 10 5 10 6 C0
port 1 nsew
rlabel  s 0 9 0 10 4 C0
port 1 nsew
rlabel  s 0 9 5 9 6 C0
port 1 nsew
rlabel  s 0 8 0 9 4 C0
port 1 nsew
rlabel  s 0 8 5 8 6 C0
port 1 nsew
rlabel  s 0 7 0 8 4 C0
port 1 nsew
rlabel  s 0 6 5 7 6 C0
port 1 nsew
rlabel  s 0 5 0 6 4 C0
port 1 nsew
rlabel  s 0 5 5 5 6 C0
port 1 nsew
rlabel  s 0 4 0 5 4 C0
port 1 nsew
rlabel  s 0 4 5 4 6 C0
port 1 nsew
rlabel  s 0 3 0 4 4 C0
port 1 nsew
rlabel  s 0 2 5 3 6 C0
port 1 nsew
rlabel  s 0 2 0 2 4 C0
port 1 nsew
rlabel  s 0 1 5 2 6 C0
port 1 nsew
rlabel  s 0 0 0 1 2 C0
port 1 nsew
rlabel  s 0 0 11 0 8 C0
port 1 nsew
rlabel  s 6 10 6 11 6 C1
port 2 nsew
rlabel  s 6 9 6 10 6 C1
port 2 nsew
rlabel  s 6 7 6 8 6 C1
port 2 nsew
rlabel  s 6 6 6 7 6 C1
port 2 nsew
rlabel  s 6 5 6 6 6 C1
port 2 nsew
rlabel  s 6 3 6 4 6 C1
port 2 nsew
rlabel  s 6 2 6 3 6 C1
port 2 nsew
rlabel  s 6 1 6 2 6 C1
port 2 nsew
rlabel  s 1 11 11 11 6 C1
port 2 nsew
rlabel  s 1 10 11 10 6 C1
port 2 nsew
rlabel  s 1 8 11 9 6 C1
port 2 nsew
rlabel  s 1 7 11 7 6 C1
port 2 nsew
rlabel  s 1 6 11 6 6 C1
port 2 nsew
rlabel  s 1 4 11 5 6 C1
port 2 nsew
rlabel  s 1 3 11 3 6 C1
port 2 nsew
rlabel  s 1 2 11 2 6 C1
port 2 nsew
rlabel  s 1 1 11 1 6 C1
port 2 nsew
rlabel r s 0 0 11 11 6 M5A
port 3 nsew
rlabel  s 0 24 0 24 4 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 11 24
string LEFview TRUE
<< end >>
