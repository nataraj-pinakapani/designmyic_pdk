magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 13 6 13 12 6 C0
port 1 nsew
rlabel  s 13 0 13 6 6 C0
port 1 nsew
rlabel  s 12 9 12 12 6 C0
port 1 nsew
rlabel  s 12 6 12 8 6 C0
port 1 nsew
rlabel  s 12 4 12 6 6 C0
port 1 nsew
rlabel  s 12 0 12 3 6 C0
port 1 nsew
rlabel  s 10 9 11 12 6 C0
port 1 nsew
rlabel  s 10 6 11 8 6 C0
port 1 nsew
rlabel  s 10 4 11 6 6 C0
port 1 nsew
rlabel  s 10 0 11 3 6 C0
port 1 nsew
rlabel  s 9 9 9 12 6 C0
port 1 nsew
rlabel  s 9 6 9 8 6 C0
port 1 nsew
rlabel  s 9 4 9 6 6 C0
port 1 nsew
rlabel  s 9 0 9 3 6 C0
port 1 nsew
rlabel  s 8 9 8 12 6 C0
port 1 nsew
rlabel  s 8 6 8 8 6 C0
port 1 nsew
rlabel  s 8 4 8 6 6 C0
port 1 nsew
rlabel  s 8 0 8 3 6 C0
port 1 nsew
rlabel  s 6 6 7 12 6 C0
port 1 nsew
rlabel  s 6 0 7 6 6 C0
port 1 nsew
rlabel  s 5 9 6 12 6 C0
port 1 nsew
rlabel  s 5 6 6 8 6 C0
port 1 nsew
rlabel  s 5 4 6 6 6 C0
port 1 nsew
rlabel  s 5 0 6 3 6 C0
port 1 nsew
rlabel  s 4 9 4 12 6 C0
port 1 nsew
rlabel  s 4 6 4 8 6 C0
port 1 nsew
rlabel  s 4 4 4 6 6 C0
port 1 nsew
rlabel  s 4 0 4 3 6 C0
port 1 nsew
rlabel  s 3 9 3 12 6 C0
port 1 nsew
rlabel  s 3 6 3 8 6 C0
port 1 nsew
rlabel  s 3 4 3 6 6 C0
port 1 nsew
rlabel  s 3 0 3 3 6 C0
port 1 nsew
rlabel  s 1 9 2 12 6 C0
port 1 nsew
rlabel  s 1 6 2 8 6 C0
port 1 nsew
rlabel  s 1 4 2 6 6 C0
port 1 nsew
rlabel  s 1 0 2 3 6 C0
port 1 nsew
rlabel  s 0 12 13 12 6 C0
port 1 nsew
rlabel  s 0 6 0 12 4 C0
port 1 nsew
rlabel  s 0 6 13 6 6 C0
port 1 nsew
rlabel  s 0 0 0 6 4 C0
port 1 nsew
rlabel  s 0 0 13 0 8 C0
port 1 nsew
rlabel  s 12 9 13 11 6 C1
port 2 nsew
rlabel  s 12 6 13 9 6 C1
port 2 nsew
rlabel  s 12 3 13 5 6 C1
port 2 nsew
rlabel  s 12 1 13 3 6 C1
port 2 nsew
rlabel  s 11 9 11 11 6 C1
port 2 nsew
rlabel  s 11 6 11 9 6 C1
port 2 nsew
rlabel  s 11 3 11 5 6 C1
port 2 nsew
rlabel  s 11 1 11 3 6 C1
port 2 nsew
rlabel  s 10 9 10 11 6 C1
port 2 nsew
rlabel  s 10 6 10 9 6 C1
port 2 nsew
rlabel  s 10 3 10 5 6 C1
port 2 nsew
rlabel  s 10 1 10 3 6 C1
port 2 nsew
rlabel  s 8 9 9 11 6 C1
port 2 nsew
rlabel  s 8 6 9 9 6 C1
port 2 nsew
rlabel  s 8 3 9 5 6 C1
port 2 nsew
rlabel  s 8 1 9 3 6 C1
port 2 nsew
rlabel  s 7 9 7 11 6 C1
port 2 nsew
rlabel  s 7 9 13 9 6 C1
port 2 nsew
rlabel  s 7 6 7 9 6 C1
port 2 nsew
rlabel  s 7 3 7 5 6 C1
port 2 nsew
rlabel  s 7 3 13 3 6 C1
port 2 nsew
rlabel  s 7 1 7 3 6 C1
port 2 nsew
rlabel  s 6 9 6 11 6 C1
port 2 nsew
rlabel  s 6 6 6 9 6 C1
port 2 nsew
rlabel  s 6 3 6 5 6 C1
port 2 nsew
rlabel  s 6 1 6 3 6 C1
port 2 nsew
rlabel  s 5 9 5 11 6 C1
port 2 nsew
rlabel  s 5 6 5 9 6 C1
port 2 nsew
rlabel  s 5 3 5 5 6 C1
port 2 nsew
rlabel  s 5 1 5 3 6 C1
port 2 nsew
rlabel  s 3 9 4 11 6 C1
port 2 nsew
rlabel  s 3 6 4 9 6 C1
port 2 nsew
rlabel  s 3 3 4 5 6 C1
port 2 nsew
rlabel  s 3 1 4 3 6 C1
port 2 nsew
rlabel  s 2 9 2 11 6 C1
port 2 nsew
rlabel  s 2 6 2 9 6 C1
port 2 nsew
rlabel  s 2 3 2 5 6 C1
port 2 nsew
rlabel  s 2 1 2 3 6 C1
port 2 nsew
rlabel  s 1 9 1 11 6 C1
port 2 nsew
rlabel  s 1 9 6 9 6 C1
port 2 nsew
rlabel  s 1 6 1 9 6 C1
port 2 nsew
rlabel  s 1 3 1 5 6 C1
port 2 nsew
rlabel  s 1 3 6 3 6 C1
port 2 nsew
rlabel  s 1 1 1 3 6 C1
port 2 nsew
rlabel  s 0 0 13 12 6 M4
port 3 nsew
rlabel metal_blue s 6 6 6 6 6 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 13 12
string LEFview TRUE
<< end >>
