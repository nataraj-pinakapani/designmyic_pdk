magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 53 75 56 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 48 75 51 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel 
 s 0 9 24 14 6 VCCD
port 3 nsew power bidirectional
rlabel 
 s 50 9 74 14 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 9 24 14 6 VCCD
port 3 nsew power bidirectional
rlabel  s 50 9 75 14 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 9 1 13 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 9 75 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 13 74 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 13 74 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 12 74 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 12 74 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 12 74 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 13 74 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 13 74 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 12 74 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 12 74 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 12 74 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 13 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 13 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 12 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 12 73 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 12 73 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 13 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 13 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 12 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 12 73 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 12 73 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 13 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 13 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 73 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 73 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 73 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 13 72 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 13 72 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 72 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 72 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 72 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 13 72 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 13 72 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 72 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 72 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 12 72 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 13 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 13 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 12 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 12 71 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 12 71 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 13 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 13 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 12 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 12 71 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 12 71 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 13 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 13 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 71 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 71 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 71 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 13 70 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 13 70 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 70 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 70 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 70 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 13 70 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 13 70 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 70 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 70 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 12 70 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 13 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 13 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 12 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 12 69 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 12 69 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 13 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 13 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 12 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 12 69 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 12 69 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 13 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 13 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 69 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 69 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 69 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 69 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 13 68 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 13 68 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 68 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 68 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 68 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 13 68 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 13 68 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 68 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 68 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 12 68 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 13 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 13 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 12 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 12 67 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 12 67 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 13 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 13 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 12 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 12 67 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 12 67 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 13 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 13 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 12 67 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 12 67 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 12 67 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 67 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 13 66 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 13 66 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 12 66 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 12 66 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 12 66 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 13 66 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 13 66 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 66 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 66 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 66 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 13 65 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 13 65 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 65 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 65 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 65 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 13 65 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 13 65 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 65 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 65 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 12 65 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 13 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 13 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 12 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 12 64 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 12 64 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 13 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 13 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 12 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 12 64 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 12 64 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 13 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 13 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 64 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 64 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 64 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 13 63 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 13 63 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 63 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 63 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 63 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 13 63 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 13 63 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 63 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 63 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 12 63 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 13 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 13 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 12 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 12 62 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 12 62 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 13 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 13 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 12 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 12 62 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 12 62 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 13 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 13 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 62 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 62 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 62 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 13 61 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 13 61 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 61 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 61 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 61 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 13 61 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 13 61 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 61 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 61 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 12 61 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 13 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 13 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 12 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 12 60 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 12 60 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 13 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 13 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 12 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 12 60 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 12 60 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 13 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 13 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 60 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 60 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 60 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 13 59 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 13 59 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 59 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 59 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 59 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 13 59 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 13 59 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 59 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 59 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 12 59 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 13 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 13 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 12 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 12 58 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 12 58 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 13 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 13 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 12 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 12 58 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 12 58 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 13 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 13 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 58 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 58 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 58 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 13 57 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 13 57 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 57 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 57 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 57 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 13 57 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 13 57 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 57 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 57 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 12 57 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 13 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 13 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 12 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 12 56 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 12 56 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 13 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 13 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 12 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 12 56 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 12 56 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 13 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 13 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 56 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 56 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 56 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 13 55 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 13 55 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 55 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 55 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 55 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 13 55 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 13 55 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 55 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 55 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 12 55 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 13 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 13 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 12 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 12 54 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 12 54 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 13 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 13 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 12 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 12 54 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 12 54 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 13 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 13 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 54 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 54 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 54 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 13 53 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 13 53 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 53 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 53 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 53 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 53 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 13 53 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 13 53 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 53 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 53 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 12 53 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 53 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 13 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 13 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 12 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 12 52 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 12 52 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 13 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 13 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 12 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 12 52 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 12 52 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 13 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 13 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 12 52 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 12 52 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 12 52 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 52 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 13 51 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 13 51 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 12 51 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 12 51 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 12 51 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 51 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 13 51 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 13 51 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 12 51 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 12 51 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 12 51 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 9 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 50 9 51 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 13 24 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 13 24 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 12 24 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 12 24 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 12 24 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 13 24 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 13 24 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 12 24 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 12 24 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 12 24 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 13 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 13 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 12 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 12 23 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 12 23 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 13 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 13 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 12 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 12 23 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 12 23 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 13 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 13 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 23 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 23 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 23 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 23 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 13 22 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 13 22 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 22 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 22 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 22 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 13 22 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 13 22 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 22 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 22 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 12 22 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 13 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 13 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 12 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 12 21 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 12 21 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 13 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 13 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 12 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 12 21 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 12 21 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 13 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 13 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 21 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 21 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 21 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 21 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 13 20 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 13 20 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 20 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 20 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 20 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 13 20 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 13 20 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 20 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 20 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 12 20 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 13 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 13 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 12 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 12 19 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 12 19 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 13 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 13 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 12 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 12 19 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 12 19 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 13 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 13 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 19 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 19 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 19 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 19 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 13 18 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 13 18 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 18 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 18 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 18 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 13 18 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 13 18 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 18 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 18 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 12 18 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 13 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 13 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 12 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 12 17 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 12 17 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 13 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 13 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 12 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 12 17 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 12 17 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 13 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 13 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 17 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 17 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 17 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 17 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 13 16 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 13 16 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 16 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 16 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 16 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 13 16 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 13 16 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 16 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 16 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 12 16 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 13 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 13 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 12 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 12 15 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 12 15 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 15 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 13 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 13 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 12 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 12 15 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 12 15 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 15 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 13 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 13 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 15 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 15 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 15 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 15 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 13 14 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 13 14 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 14 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 14 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 14 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 13 14 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 13 14 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 14 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 14 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 12 14 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 13 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 13 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 12 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 12 13 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 12 13 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 13 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 13 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 12 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 12 13 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 12 13 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 13 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 13 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 13 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 13 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 13 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 13 12 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 13 12 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 12 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 12 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 12 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 13 12 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 13 12 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 12 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 12 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 12 12 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 13 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 13 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 12 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 12 11 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 12 11 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 13 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 13 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 12 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 12 11 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 12 11 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 13 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 13 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 11 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 11 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 11 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 13 10 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 13 10 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 10 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 10 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 10 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 13 10 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 13 10 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 10 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 10 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 12 10 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 13 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 13 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 12 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 12 9 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 12 9 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 13 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 13 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 12 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 12 9 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 12 9 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 13 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 13 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 9 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 9 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 9 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 13 8 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 13 8 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 8 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 8 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 8 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 13 8 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 13 8 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 8 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 8 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 12 8 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 13 7 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 13 7 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 12 7 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 12 7 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 12 7 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 13 7 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 13 7 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 12 7 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 12 7 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 12 7 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 13 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 13 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 12 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 12 6 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 12 6 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 13 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 13 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 12 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 12 6 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 12 6 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 13 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 13 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 6 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 6 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 6 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 6 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 13 5 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 13 5 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 5 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 5 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 5 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 13 5 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 13 5 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 5 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 5 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 12 5 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 13 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 13 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 12 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 12 4 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 12 4 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 13 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 13 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 12 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 12 4 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 12 4 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 13 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 13 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 4 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 4 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 4 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 4 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 13 3 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 13 3 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 3 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 3 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 3 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 13 3 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 13 3 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 3 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 3 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 12 3 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 13 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 13 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 12 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 12 2 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 12 2 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 13 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 13 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 12 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 12 2 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 12 2 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 13 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 13 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 2 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 2 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 2 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 2 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 13 1 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 13 1 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 1 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 1 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 1 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 13 1 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 13 1 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 1 13 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 1 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 12 1 12 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 9 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 69 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 64 1 68 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 68 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 1 48 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 52 1 53 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 56 1 57 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 48 75 48 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 52 75 53 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 56 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 1 57 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 48 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
