/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1.spice