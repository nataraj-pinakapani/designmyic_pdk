magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 10 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 10 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 46 10 55 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 54 10 55 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 46 10 46 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 35 10 38 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 35 10 38 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 13 10 16 6 VDDA
port 4 nsew power bidirectional
rlabel  s 0 13 10 16 6 VDDA
port 4 nsew power bidirectional
rlabel  s 0 30 10 33 6 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 30 10 33 6 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 62 10 66 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 62 10 67 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 0 10 5 6 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 0 10 5 6 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 68 10 93 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 68 10 93 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 18 10 22 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 18 10 22 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 7 10 11 6 VCCD
port 9 nsew power bidirectional
rlabel  s 0 7 10 12 6 VCCD
port 9 nsew power bidirectional
rlabel  s 0 24 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 10 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 10 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 40 10 44 6 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 40 10 44 6 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 56 10 61 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 56 10 61 6 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string LEFclass PAD SPACER
string FIXED_BBOX 0 0 10 198
string LEFview TRUE
<< end >>
