magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 39 21 582 157
rect 39 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 125 47 155 131
rect 211 47 241 131
rect 311 47 341 131
rect 397 47 427 131
rect 469 47 499 131
<< scpmoshvt >>
rect 139 369 169 497
rect 211 369 241 497
rect 283 369 313 497
rect 369 369 399 497
rect 475 369 505 497
<< ndiff >>
rect 65 93 125 131
rect 65 59 73 93
rect 107 59 125 93
rect 65 47 125 59
rect 155 101 211 131
rect 155 67 166 101
rect 200 67 211 101
rect 155 47 211 67
rect 241 89 311 131
rect 241 55 258 89
rect 292 55 311 89
rect 241 47 311 55
rect 341 106 397 131
rect 341 72 352 106
rect 386 72 397 106
rect 341 47 397 72
rect 427 47 469 131
rect 499 89 556 131
rect 499 55 510 89
rect 544 55 556 89
rect 499 47 556 55
<< pdiff >>
rect 80 483 139 497
rect 80 449 88 483
rect 122 449 139 483
rect 80 415 139 449
rect 80 381 88 415
rect 122 381 139 415
rect 80 369 139 381
rect 169 369 211 497
rect 241 369 283 497
rect 313 483 369 497
rect 313 449 324 483
rect 358 449 369 483
rect 313 415 369 449
rect 313 381 324 415
rect 358 381 369 415
rect 313 369 369 381
rect 399 485 475 497
rect 399 451 424 485
rect 458 451 475 485
rect 399 369 475 451
rect 505 483 566 497
rect 505 449 524 483
rect 558 449 566 483
rect 505 415 566 449
rect 505 381 524 415
rect 558 381 566 415
rect 505 369 566 381
<< ndiffc >>
rect 73 59 107 93
rect 166 67 200 101
rect 258 55 292 89
rect 352 72 386 106
rect 510 55 544 89
<< pdiffc >>
rect 88 449 122 483
rect 88 381 122 415
rect 324 449 358 483
rect 324 381 358 415
rect 424 451 458 485
rect 524 449 558 483
rect 524 381 558 415
<< poly >>
rect 139 497 169 523
rect 211 497 241 523
rect 283 497 313 523
rect 369 497 399 523
rect 475 497 505 523
rect 139 354 169 369
rect 43 324 169 354
rect 43 280 97 324
rect 211 282 241 369
rect 43 246 53 280
rect 87 246 97 280
rect 43 203 97 246
rect 175 261 241 282
rect 175 227 191 261
rect 225 227 241 261
rect 175 213 241 227
rect 43 169 53 203
rect 87 176 97 203
rect 87 169 155 176
rect 43 146 155 169
rect 125 131 155 146
rect 211 131 241 213
rect 283 279 313 369
rect 369 354 399 369
rect 475 354 505 369
rect 369 319 433 354
rect 475 324 623 354
rect 395 282 433 319
rect 567 316 623 324
rect 567 282 579 316
rect 613 282 623 316
rect 283 261 353 279
rect 283 227 305 261
rect 339 227 353 261
rect 283 211 353 227
rect 395 264 525 282
rect 395 230 407 264
rect 441 230 475 264
rect 509 230 525 264
rect 395 218 525 230
rect 567 248 623 282
rect 395 211 427 218
rect 311 131 341 211
rect 397 131 427 211
rect 567 214 579 248
rect 613 214 623 248
rect 567 176 623 214
rect 469 146 623 176
rect 469 131 499 146
rect 125 21 155 47
rect 211 21 241 47
rect 311 21 341 47
rect 397 21 427 47
rect 469 21 499 47
<< polycont >>
rect 53 246 87 280
rect 191 227 225 261
rect 53 169 87 203
rect 579 282 613 316
rect 305 227 339 261
rect 407 230 441 264
rect 475 230 509 264
rect 579 214 613 248
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 72 483 157 493
rect 72 449 88 483
rect 122 449 157 483
rect 308 483 374 493
rect 72 415 157 449
rect 72 381 88 415
rect 122 381 157 415
rect 72 365 157 381
rect 17 280 87 331
rect 17 246 53 280
rect 17 203 87 246
rect 17 169 53 203
rect 17 146 87 169
rect 121 177 157 365
rect 191 261 265 472
rect 308 449 324 483
rect 358 449 374 483
rect 408 485 474 527
rect 408 451 424 485
rect 458 451 474 485
rect 508 483 574 493
rect 308 417 374 449
rect 508 449 524 483
rect 558 449 574 483
rect 508 417 574 449
rect 308 415 574 417
rect 308 381 324 415
rect 358 381 524 415
rect 558 381 574 415
rect 225 227 265 261
rect 191 211 265 227
rect 299 261 369 347
rect 471 280 525 347
rect 299 227 305 261
rect 339 227 369 261
rect 299 211 369 227
rect 407 264 525 280
rect 441 230 475 264
rect 509 230 525 264
rect 407 214 525 230
rect 121 127 408 177
rect 471 132 525 214
rect 559 316 627 347
rect 559 282 579 316
rect 613 282 627 316
rect 559 248 627 282
rect 559 214 579 248
rect 613 214 627 248
rect 559 130 627 214
rect 157 123 408 127
rect 157 101 208 123
rect 57 59 73 93
rect 107 59 123 93
rect 57 17 123 59
rect 157 67 166 101
rect 200 67 208 101
rect 342 106 408 123
rect 157 51 208 67
rect 242 55 258 89
rect 292 55 308 89
rect 342 72 352 106
rect 386 72 408 106
rect 342 56 408 72
rect 494 89 560 96
rect 242 17 308 55
rect 494 55 510 89
rect 544 55 560 89
rect 494 17 560 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 581 153 615 187 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 121 425 155 459 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 121 357 155 391 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 121 289 155 323 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 121 221 155 255 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 121 153 155 187 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 213 289 247 323 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 213 357 247 391 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 213 425 247 459 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 489 153 523 187 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 a2111oi_0
rlabel metal1 s 0 -48 644 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3790586
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3783122
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 16.100 13.600 
<< end >>
