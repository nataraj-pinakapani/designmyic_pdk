magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 9 -205 12 -202 8 B_P
port 1 nsew
rlabel  s 105 102 109 103 6 D_N2
port 2 nsew
rlabel  s 104 102 104 103 6 D_N2
port 2 nsew
rlabel  s 103 102 104 103 6 D_N2
port 2 nsew
rlabel  s 102 103 109 103 6 D_N2
port 2 nsew
rlabel  s 102 102 103 103 6 D_N2
port 2 nsew
rlabel  s 68 -125 69 -125 8 D_P
port 3 nsew
rlabel  s 101 -123 103 -122 8 D_P2
port 4 nsew
rlabel  s 69 100 70 101 6 G
port 5 nsew
rlabel  s 102 103 105 112 6 G_N2
port 6 nsew
rlabel  s 68 -124 69 -124 8 G_P
port 7 nsew
rlabel  s 103 -122 104 -121 8 G_P2
port 8 nsew
rlabel  s 9 9 12 12 6 NWELL
port 9 nsew
rlabel  s 70 100 70 100 6 S
port 10 nsew
rlabel  s 69 100 69 100 6 S
port 10 nsew
rlabel  s 69 99 70 100 6 S
port 10 nsew
rlabel  s 105 100 106 103 6 S_N2
port 11 nsew
rlabel  s 105 100 105 103 6 S_N2
port 11 nsew
rlabel  s 104 100 104 103 6 S_N2
port 11 nsew
rlabel  s 103 100 103 103 6 S_N2
port 11 nsew
rlabel  s 102 100 102 103 6 S_N2
port 11 nsew
rlabel  s 102 88 106 100 6 S_N2
port 11 nsew
rlabel  s 69 -126 69 -125 8 S_P
port 12 nsew
rlabel  s 68 -126 68 -125 8 S_P
port 12 nsew
rlabel  s 68 -126 69 -126 8 S_P
port 12 nsew
rlabel  s 104 -126 104 -122 8 S_P2
port 13 nsew
rlabel  s 103 -126 103 -122 8 S_P2
port 13 nsew
rlabel  s 103 -127 104 -126 8 S_P2
port 13 nsew
rlabel  s 60 91 63 94 6 VGND
port 14 nsew ground default
rlabel  s 69 100 70 100 6 VPWR
port 15 nsew power default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 -214 1556 198
string LEFview TRUE
<< end >>
