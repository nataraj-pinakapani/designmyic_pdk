magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 34 201 1433 203
rect 34 23 1744 201
rect 34 21 247 23
rect 744 21 936 23
rect 1348 21 1744 23
rect 34 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 112 47 142 177
rect 236 93 266 177
rect 458 49 488 177
rect 568 49 598 177
rect 830 47 860 177
rect 1016 49 1046 177
rect 1168 49 1198 133
rect 1327 49 1357 177
rect 1447 47 1477 167
rect 1547 47 1577 175
rect 1631 47 1661 175
<< scpmoshvt >>
rect 116 297 146 497
rect 236 297 266 425
rect 450 325 480 493
rect 556 325 586 493
rect 797 297 827 497
rect 1016 297 1046 465
rect 1168 297 1198 425
rect 1343 329 1373 457
rect 1446 329 1476 497
rect 1547 297 1577 497
rect 1631 297 1661 497
<< ndiff >>
rect 60 129 112 177
rect 60 95 68 129
rect 102 95 112 129
rect 60 47 112 95
rect 142 93 236 177
rect 266 169 350 177
rect 266 135 304 169
rect 338 135 350 169
rect 266 93 350 135
rect 404 165 458 177
rect 404 131 414 165
rect 448 131 458 165
rect 142 89 221 93
rect 142 55 168 89
rect 202 55 221 89
rect 142 47 221 55
rect 404 49 458 131
rect 488 91 568 177
rect 488 57 498 91
rect 532 57 568 91
rect 488 49 568 57
rect 598 169 697 177
rect 598 135 650 169
rect 684 135 697 169
rect 598 49 697 135
rect 770 157 830 177
rect 770 123 786 157
rect 820 123 830 157
rect 770 89 830 123
rect 770 55 786 89
rect 820 55 830 89
rect 770 47 830 55
rect 860 161 912 177
rect 860 127 870 161
rect 904 127 912 161
rect 860 121 912 127
rect 860 47 910 121
rect 966 105 1016 177
rect 964 97 1016 105
rect 964 63 972 97
rect 1006 63 1016 97
rect 964 49 1016 63
rect 1046 133 1147 177
rect 1223 169 1327 177
rect 1223 135 1269 169
rect 1303 135 1327 169
rect 1223 133 1327 135
rect 1046 126 1168 133
rect 1046 92 1056 126
rect 1090 92 1168 126
rect 1046 49 1168 92
rect 1198 49 1327 133
rect 1357 167 1407 177
rect 1497 167 1547 175
rect 1357 93 1447 167
rect 1357 59 1369 93
rect 1403 59 1447 93
rect 1357 49 1447 59
rect 1374 47 1447 49
rect 1477 142 1547 167
rect 1477 108 1503 142
rect 1537 108 1547 142
rect 1477 47 1547 108
rect 1577 97 1631 175
rect 1577 63 1587 97
rect 1621 63 1631 97
rect 1577 47 1631 63
rect 1661 101 1718 175
rect 1661 67 1671 101
rect 1705 67 1718 101
rect 1661 47 1718 67
<< pdiff >>
rect 60 477 116 497
rect 60 443 72 477
rect 106 443 116 477
rect 60 409 116 443
rect 60 375 72 409
rect 106 375 116 409
rect 60 341 116 375
rect 60 307 72 341
rect 106 307 116 341
rect 60 297 116 307
rect 146 477 221 497
rect 146 443 173 477
rect 207 443 221 477
rect 146 425 221 443
rect 146 297 236 425
rect 266 341 322 425
rect 266 307 276 341
rect 310 307 322 341
rect 386 413 450 493
rect 386 379 406 413
rect 440 379 450 413
rect 386 325 450 379
rect 480 481 556 493
rect 480 447 499 481
rect 533 447 556 481
rect 480 325 556 447
rect 586 481 691 493
rect 586 447 646 481
rect 680 447 691 481
rect 586 325 691 447
rect 745 481 797 497
rect 745 447 753 481
rect 787 447 797 481
rect 266 297 322 307
rect 745 297 797 447
rect 827 349 877 497
rect 931 405 1016 465
rect 931 371 939 405
rect 973 371 1016 405
rect 931 365 1016 371
rect 827 343 879 349
rect 827 309 837 343
rect 871 309 879 343
rect 827 297 879 309
rect 933 297 1016 365
rect 1046 425 1146 465
rect 1388 489 1446 497
rect 1388 457 1400 489
rect 1258 425 1343 457
rect 1046 409 1168 425
rect 1046 375 1097 409
rect 1131 375 1168 409
rect 1046 341 1168 375
rect 1046 307 1097 341
rect 1131 307 1168 341
rect 1046 297 1168 307
rect 1198 421 1343 425
rect 1198 387 1299 421
rect 1333 387 1343 421
rect 1198 329 1343 387
rect 1373 455 1400 457
rect 1434 455 1446 489
rect 1373 329 1446 455
rect 1476 341 1547 497
rect 1476 329 1503 341
rect 1198 297 1293 329
rect 1491 307 1503 329
rect 1537 307 1547 341
rect 1491 297 1547 307
rect 1577 489 1631 497
rect 1577 455 1587 489
rect 1621 455 1631 489
rect 1577 297 1631 455
rect 1661 477 1718 497
rect 1661 443 1672 477
rect 1706 443 1718 477
rect 1661 409 1718 443
rect 1661 375 1672 409
rect 1706 375 1718 409
rect 1661 297 1718 375
<< ndiffc >>
rect 68 95 102 129
rect 304 135 338 169
rect 414 131 448 165
rect 168 55 202 89
rect 498 57 532 91
rect 650 135 684 169
rect 786 123 820 157
rect 786 55 820 89
rect 870 127 904 161
rect 972 63 1006 97
rect 1269 135 1303 169
rect 1056 92 1090 126
rect 1369 59 1403 93
rect 1503 108 1537 142
rect 1587 63 1621 97
rect 1671 67 1705 101
<< pdiffc >>
rect 72 443 106 477
rect 72 375 106 409
rect 72 307 106 341
rect 173 443 207 477
rect 276 307 310 341
rect 406 379 440 413
rect 499 447 533 481
rect 646 447 680 481
rect 753 447 787 481
rect 939 371 973 405
rect 837 309 871 343
rect 1097 375 1131 409
rect 1097 307 1131 341
rect 1299 387 1333 421
rect 1400 455 1434 489
rect 1503 307 1537 341
rect 1587 455 1621 489
rect 1672 443 1706 477
rect 1672 375 1706 409
<< poly >>
rect 116 497 146 523
rect 450 493 480 519
rect 556 493 586 519
rect 797 497 827 523
rect 236 425 266 483
rect 116 265 146 297
rect 236 265 266 297
rect 450 271 480 325
rect 450 265 489 271
rect 556 265 586 325
rect 1016 493 1373 523
rect 1446 497 1476 523
rect 1547 497 1577 523
rect 1631 497 1661 523
rect 1016 465 1046 493
rect 1343 457 1373 493
rect 1168 425 1198 451
rect 112 249 194 265
rect 112 215 150 249
rect 184 215 194 249
rect 112 199 194 215
rect 236 249 489 265
rect 236 215 377 249
rect 411 215 445 249
rect 479 215 489 249
rect 236 199 489 215
rect 544 249 598 265
rect 544 215 554 249
rect 588 215 598 249
rect 797 247 827 297
rect 1016 247 1046 297
rect 1168 265 1198 297
rect 1343 265 1373 329
rect 797 217 1046 247
rect 544 199 598 215
rect 112 177 142 199
rect 236 177 266 199
rect 458 197 489 199
rect 458 177 488 197
rect 568 177 598 199
rect 830 177 860 217
rect 1016 177 1046 217
rect 1088 249 1198 265
rect 1088 215 1098 249
rect 1132 215 1198 249
rect 1088 199 1198 215
rect 236 67 266 93
rect 112 21 142 47
rect 458 21 488 49
rect 568 21 598 49
rect 1168 133 1198 199
rect 1327 249 1381 265
rect 1446 256 1476 329
rect 1547 265 1577 297
rect 1631 265 1661 297
rect 1446 255 1477 256
rect 1327 215 1337 249
rect 1371 215 1381 249
rect 1327 199 1381 215
rect 1423 239 1477 255
rect 1423 205 1433 239
rect 1467 205 1477 239
rect 1327 177 1357 199
rect 1423 189 1477 205
rect 1519 249 1577 265
rect 1519 215 1529 249
rect 1563 215 1577 249
rect 1519 199 1577 215
rect 1619 249 1673 265
rect 1619 215 1629 249
rect 1663 215 1673 249
rect 1619 199 1673 215
rect 1447 167 1477 189
rect 1547 175 1577 199
rect 1631 175 1661 199
rect 830 21 860 47
rect 1016 21 1046 49
rect 1168 23 1198 49
rect 1327 21 1357 49
rect 1447 21 1477 47
rect 1547 21 1577 47
rect 1631 21 1661 47
<< polycont >>
rect 150 215 184 249
rect 377 215 411 249
rect 445 215 479 249
rect 554 215 588 249
rect 1098 215 1132 249
rect 1337 215 1371 249
rect 1433 205 1467 239
rect 1529 215 1563 249
rect 1629 215 1663 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 17 477 122 493
rect 17 443 72 477
rect 106 443 122 477
rect 156 477 223 527
rect 737 481 803 527
rect 1571 489 1638 527
rect 156 443 173 477
rect 207 443 223 477
rect 260 447 499 481
rect 533 447 579 481
rect 622 447 646 481
rect 680 447 703 481
rect 737 447 753 481
rect 787 447 803 481
rect 870 455 1400 489
rect 1434 455 1489 489
rect 1571 455 1587 489
rect 1621 455 1638 489
rect 1672 477 1731 493
rect 17 409 122 443
rect 260 409 294 447
rect 669 413 703 447
rect 870 413 904 455
rect 17 375 72 409
rect 106 375 122 409
rect 17 341 122 375
rect 17 307 72 341
rect 106 307 122 341
rect 17 288 122 307
rect 156 375 294 409
rect 374 379 406 413
rect 440 379 635 413
rect 669 379 904 413
rect 939 405 973 421
rect 17 185 80 288
rect 156 265 190 375
rect 237 307 276 341
rect 310 307 567 341
rect 150 249 190 265
rect 184 215 190 249
rect 150 199 190 215
rect 17 129 118 185
rect 156 173 190 199
rect 156 139 270 173
rect 17 95 68 129
rect 102 95 118 129
rect 17 70 118 95
rect 152 89 202 105
rect 152 55 168 89
rect 152 17 202 55
rect 236 85 270 139
rect 304 169 338 307
rect 533 265 567 307
rect 601 339 635 379
rect 601 323 707 339
rect 601 305 673 323
rect 650 289 673 305
rect 650 275 707 289
rect 372 249 499 265
rect 372 215 377 249
rect 411 215 445 249
rect 479 215 499 249
rect 372 199 499 215
rect 533 249 588 265
rect 533 215 554 249
rect 533 199 588 215
rect 650 169 684 275
rect 741 241 775 379
rect 821 309 837 343
rect 871 309 904 343
rect 821 289 904 309
rect 304 119 338 135
rect 394 131 414 165
rect 448 131 616 165
rect 478 85 498 91
rect 236 57 498 85
rect 532 57 548 91
rect 236 51 548 57
rect 582 85 616 131
rect 650 119 684 135
rect 718 207 775 241
rect 718 85 752 207
rect 856 187 904 289
rect 582 51 752 85
rect 786 157 820 173
rect 786 89 820 123
rect 856 153 857 187
rect 891 161 904 187
rect 856 127 870 153
rect 856 83 904 127
rect 939 119 973 371
rect 1007 178 1041 455
rect 1706 443 1731 477
rect 1672 421 1731 443
rect 1079 375 1097 409
rect 1131 375 1162 409
rect 1079 341 1162 375
rect 1079 307 1097 341
rect 1131 323 1162 341
rect 1269 387 1299 421
rect 1333 409 1731 421
rect 1333 387 1672 409
rect 1131 307 1133 323
rect 1079 289 1133 307
rect 1167 289 1235 323
rect 1082 249 1167 254
rect 1082 215 1098 249
rect 1132 215 1167 249
rect 1082 199 1167 215
rect 1124 187 1167 199
rect 1007 165 1051 178
rect 1007 144 1090 165
rect 1017 131 1090 144
rect 1056 126 1090 131
rect 1124 153 1133 187
rect 1124 126 1167 153
rect 939 85 949 119
rect 786 17 820 55
rect 939 63 972 85
rect 1006 63 1022 97
rect 1056 64 1090 92
rect 1201 85 1235 289
rect 1269 169 1303 387
rect 1634 375 1672 387
rect 1706 375 1731 409
rect 1337 289 1453 323
rect 1487 307 1503 341
rect 1537 307 1651 341
rect 1487 299 1651 307
rect 1337 249 1371 289
rect 1617 265 1651 299
rect 1337 199 1371 215
rect 1405 239 1467 255
rect 1405 205 1433 239
rect 1501 249 1583 265
rect 1501 215 1529 249
rect 1563 215 1583 249
rect 1617 249 1663 265
rect 1617 215 1629 249
rect 1405 189 1467 205
rect 1617 199 1663 215
rect 1405 187 1446 189
rect 1405 153 1409 187
rect 1443 153 1446 187
rect 1617 181 1651 199
rect 1405 146 1446 153
rect 1503 150 1651 181
rect 1495 147 1651 150
rect 1269 119 1303 135
rect 1495 142 1553 147
rect 1495 119 1503 142
rect 1337 85 1369 93
rect 939 53 1022 63
rect 1201 59 1369 85
rect 1403 59 1430 93
rect 1495 85 1501 119
rect 1537 108 1553 142
rect 1697 117 1731 375
rect 1535 85 1553 108
rect 1495 59 1553 85
rect 1587 97 1621 113
rect 1201 51 1430 59
rect 1587 17 1621 63
rect 1671 101 1731 117
rect 1705 67 1731 101
rect 1671 51 1731 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 673 289 707 323
rect 857 161 891 187
rect 857 153 870 161
rect 870 153 891 161
rect 1133 289 1167 323
rect 1133 153 1167 187
rect 949 97 983 119
rect 949 85 972 97
rect 972 85 983 97
rect 1409 153 1443 187
rect 1501 108 1503 119
rect 1503 108 1535 119
rect 1501 85 1535 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 661 323 719 329
rect 661 289 673 323
rect 707 320 719 323
rect 1121 323 1179 329
rect 1121 320 1133 323
rect 707 292 1133 320
rect 707 289 719 292
rect 661 283 719 289
rect 1121 289 1133 292
rect 1167 289 1179 323
rect 1121 283 1179 289
rect 845 187 903 193
rect 845 153 857 187
rect 891 184 903 187
rect 1121 187 1179 193
rect 1121 184 1133 187
rect 891 156 1133 184
rect 891 153 903 156
rect 845 147 903 153
rect 1121 153 1133 156
rect 1167 184 1179 187
rect 1397 187 1455 193
rect 1397 184 1409 187
rect 1167 156 1409 184
rect 1167 153 1179 156
rect 1121 147 1179 153
rect 1397 153 1409 156
rect 1443 153 1455 187
rect 1397 147 1455 153
rect 937 119 995 125
rect 937 85 949 119
rect 983 116 995 119
rect 1489 119 1547 125
rect 1489 116 1501 119
rect 983 88 1501 116
rect 983 85 995 88
rect 937 79 995 85
rect 1489 85 1501 88
rect 1535 85 1547 119
rect 1489 79 1547 85
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1409 289 1443 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1501 221 1535 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 xor3_1
rlabel metal1 s 0 -48 1748 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_END 673232
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 661420
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 8.740 0.000 
<< end >>
