magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 4 3 6 6 DRAIN
port 1 nsew
rlabel rotate s 2 7 2 7 6 GATE
port 2 nsew
rlabel rotate s 2 6 2 6 6 GATE
port 2 nsew
rlabel rotate s 2 0 2 1 8 GATE
port 2 nsew
rlabel rotate s 2 0 2 0 8 GATE
port 2 nsew
rlabel rotate s 1 7 2 7 6 GATE
port 2 nsew
rlabel rotate s 1 6 2 6 6 GATE
port 2 nsew
rlabel rotate s 1 0 2 1 8 GATE
port 2 nsew
rlabel rotate s 1 0 2 0 8 GATE
port 2 nsew
rlabel  s 1 6 2 7 6 GATE
port 2 nsew
rlabel  s 1 0 2 1 8 GATE
port 2 nsew
rlabel  s 1 6 2 7 6 GATE
port 2 nsew
rlabel  s 1 0 2 1 8 GATE
port 2 nsew
rlabel  s 0 1 3 3 6 SOURCE
port 3 nsew
rlabel  s 0 1 1 6 4 SUBSTRATE
port 4 nsew
rlabel  s 3 1 3 6 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 3 7
string LEFview TRUE
<< end >>
