/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/fixed_devices/sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50_fail.cdl