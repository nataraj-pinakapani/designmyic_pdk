magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< pwell >>
rect 0 643 796 796
rect 0 153 153 643
rect 643 153 796 643
rect 0 0 796 153
<< nbase >>
rect 153 153 643 643
<< pdiff >>
rect 330 449 466 466
rect 330 347 347 449
rect 449 347 466 449
rect 330 330 466 347
<< pdiffc >>
rect 347 347 449 449
<< psubdiff >>
rect 26 736 770 770
rect 26 702 60 736
rect 94 702 128 736
rect 162 702 196 736
rect 230 702 264 736
rect 298 702 498 736
rect 532 702 566 736
rect 600 702 634 736
rect 668 702 702 736
rect 736 702 770 736
rect 26 669 770 702
rect 26 668 127 669
rect 26 634 60 668
rect 94 634 127 668
rect 26 600 127 634
rect 669 668 770 669
rect 669 634 702 668
rect 736 634 770 668
rect 26 566 60 600
rect 94 566 127 600
rect 26 532 127 566
rect 26 498 60 532
rect 94 498 127 532
rect 26 298 127 498
rect 26 264 60 298
rect 94 264 127 298
rect 26 230 127 264
rect 26 196 60 230
rect 94 196 127 230
rect 26 162 127 196
rect 669 600 770 634
rect 669 566 702 600
rect 736 566 770 600
rect 669 532 770 566
rect 669 498 702 532
rect 736 498 770 532
rect 669 298 770 498
rect 669 264 702 298
rect 736 264 770 298
rect 669 230 770 264
rect 669 196 702 230
rect 736 196 770 230
rect 26 128 60 162
rect 94 128 127 162
rect 26 127 127 128
rect 669 162 770 196
rect 669 128 702 162
rect 736 128 770 162
rect 669 127 770 128
rect 26 94 770 127
rect 26 60 60 94
rect 94 60 128 94
rect 162 60 196 94
rect 230 60 264 94
rect 298 60 498 94
rect 532 60 566 94
rect 600 60 634 94
rect 668 60 702 94
rect 736 60 770 94
rect 26 26 770 60
<< nsubdiff >>
rect 189 583 607 607
rect 189 549 213 583
rect 247 549 281 583
rect 315 549 481 583
rect 515 549 549 583
rect 583 549 607 583
rect 189 535 607 549
rect 189 515 261 535
rect 189 481 213 515
rect 247 481 261 515
rect 189 315 261 481
rect 535 515 607 535
rect 535 481 549 515
rect 583 481 607 515
rect 189 281 213 315
rect 247 281 261 315
rect 189 261 261 281
rect 535 315 607 481
rect 535 281 549 315
rect 583 281 607 315
rect 535 261 607 281
rect 189 247 607 261
rect 189 213 213 247
rect 247 213 281 247
rect 315 213 481 247
rect 515 213 549 247
rect 583 213 607 247
rect 189 189 607 213
<< psubdiffcont >>
rect 60 702 94 736
rect 128 702 162 736
rect 196 702 230 736
rect 264 702 298 736
rect 498 702 532 736
rect 566 702 600 736
rect 634 702 668 736
rect 702 702 736 736
rect 60 634 94 668
rect 702 634 736 668
rect 60 566 94 600
rect 60 498 94 532
rect 60 264 94 298
rect 60 196 94 230
rect 702 566 736 600
rect 702 498 736 532
rect 702 264 736 298
rect 702 196 736 230
rect 60 128 94 162
rect 702 128 736 162
rect 60 60 94 94
rect 128 60 162 94
rect 196 60 230 94
rect 264 60 298 94
rect 498 60 532 94
rect 566 60 600 94
rect 634 60 668 94
rect 702 60 736 94
<< nsubdiffcont >>
rect 213 549 247 583
rect 281 549 315 583
rect 481 549 515 583
rect 549 549 583 583
rect 213 481 247 515
rect 549 481 583 515
rect 213 281 247 315
rect 549 281 583 315
rect 213 213 247 247
rect 281 213 315 247
rect 481 213 515 247
rect 549 213 583 247
<< locali >>
rect 26 736 770 770
rect 26 702 60 736
rect 94 702 128 736
rect 162 702 196 736
rect 230 702 264 736
rect 298 702 498 736
rect 532 702 566 736
rect 600 702 634 736
rect 668 702 702 736
rect 736 702 770 736
rect 26 669 770 702
rect 26 668 127 669
rect 26 634 60 668
rect 94 634 127 668
rect 26 600 127 634
rect 669 668 770 669
rect 669 634 702 668
rect 736 634 770 668
rect 26 566 60 600
rect 94 566 127 600
rect 26 532 127 566
rect 26 498 60 532
rect 94 498 127 532
rect 26 298 127 498
rect 26 264 60 298
rect 94 264 127 298
rect 26 230 127 264
rect 26 196 60 230
rect 94 196 127 230
rect 26 162 127 196
rect 189 583 607 607
rect 189 549 213 583
rect 247 549 281 583
rect 315 549 481 583
rect 515 549 549 583
rect 583 549 607 583
rect 189 535 607 549
rect 189 515 261 535
rect 189 481 213 515
rect 247 481 261 515
rect 189 315 261 481
rect 535 515 607 535
rect 535 481 549 515
rect 583 481 607 515
rect 319 463 477 477
rect 319 429 333 463
rect 367 449 429 463
rect 463 429 477 463
rect 319 367 347 429
rect 449 367 477 429
rect 319 333 333 367
rect 367 333 429 347
rect 463 333 477 367
rect 319 319 477 333
rect 189 281 213 315
rect 247 281 261 315
rect 189 261 261 281
rect 535 315 607 481
rect 535 281 549 315
rect 583 281 607 315
rect 535 261 607 281
rect 189 247 607 261
rect 189 213 213 247
rect 247 213 281 247
rect 315 213 481 247
rect 515 213 549 247
rect 583 213 607 247
rect 189 189 607 213
rect 669 600 770 634
rect 669 566 702 600
rect 736 566 770 600
rect 669 532 770 566
rect 669 498 702 532
rect 736 498 770 532
rect 669 298 770 498
rect 669 264 702 298
rect 736 264 770 298
rect 669 230 770 264
rect 669 196 702 230
rect 736 196 770 230
rect 26 128 60 162
rect 94 128 127 162
rect 26 127 127 128
rect 669 162 770 196
rect 669 128 702 162
rect 736 128 770 162
rect 669 127 770 128
rect 26 94 770 127
rect 26 60 60 94
rect 94 60 128 94
rect 162 60 196 94
rect 230 60 264 94
rect 298 60 498 94
rect 532 60 566 94
rect 600 60 634 94
rect 668 60 702 94
rect 736 60 770 94
rect 26 26 770 60
<< viali >>
rect 333 449 367 463
rect 429 449 463 463
rect 333 429 347 449
rect 347 429 367 449
rect 429 429 449 449
rect 449 429 463 449
rect 333 347 347 367
rect 347 347 367 367
rect 429 347 449 367
rect 449 347 463 367
rect 333 333 367 347
rect 429 333 463 347
<< metal1 >>
rect 315 463 481 481
rect 315 429 333 463
rect 367 429 429 463
rect 463 429 481 463
rect 315 367 481 429
rect 315 333 333 367
rect 367 333 429 367
rect 463 333 481 367
rect 315 315 481 333
<< comment >>
rect 26 782 27 795
tri 27 782 31 786 se
tri 765 782 769 786 sw
rect 769 782 770 795
rect 26 781 371 782
rect 424 781 770 782
rect 26 769 27 781
tri 27 777 31 781 ne
tri 765 777 769 781 nw
rect 769 769 770 781
rect 153 620 154 633
tri 154 620 158 624 se
tri 638 620 642 624 sw
rect 642 620 643 633
rect 153 619 345 620
rect 452 619 643 620
rect 153 607 154 619
tri 154 615 158 619 ne
tri 638 615 642 619 nw
rect 642 607 643 619
rect 189 565 190 578
tri 190 565 194 569 se
tri 208 565 212 569 sw
rect 212 565 213 578
rect 189 564 213 565
rect 189 552 190 564
tri 190 560 194 564 ne
rect 208 563 211 564
tri 211 563 212 564 nw
tri 199 560 201 563 se
tri 208 560 211 563 nw
tri 198 557 199 560 se
rect 199 557 201 560
tri 201 557 202 560 sw
rect 197 556 198 557
tri 198 556 199 557 nw
rect 201 556 202 557
rect 195 524 200 556
rect 212 552 213 564
rect 607 533 608 546
tri 608 533 612 537 se
tri 664 533 668 537 sw
rect 668 533 669 546
rect 607 532 669 533
rect 607 520 608 532
tri 608 528 612 532 ne
tri 664 528 668 532 nw
rect 668 520 669 532
rect 330 479 331 492
tri 331 479 335 483 se
tri 461 479 465 483 sw
rect 465 479 466 492
rect 330 478 377 479
rect 419 478 466 479
rect 330 466 331 478
tri 331 474 335 478 ne
tri 461 474 465 478 nw
rect 465 466 466 478
rect 189 442 190 455
tri 190 442 194 446 se
tri 256 442 260 446 sw
rect 260 442 261 455
rect 189 441 261 442
rect 189 429 190 441
tri 190 437 194 441 ne
tri 256 437 260 441 nw
rect 260 429 261 441
tri 390 404 392 406 se
tri 392 404 393 406 sw
tri 403 404 404 406 se
tri 404 404 406 406 sw
tri 390 403 392 404 ne
rect 392 403 393 404
tri 393 403 395 404 sw
tri 401 403 403 404 se
tri 392 400 395 403 ne
tri 395 401 396 403 sw
tri 400 401 401 403 se
rect 401 401 403 403
tri 403 401 406 404 nw
rect 395 400 396 401
tri 396 400 398 401 sw
tri 398 400 400 401 se
tri 395 398 396 400 ne
tri 393 395 396 398 se
rect 396 396 400 400
tri 400 398 403 401 nw
rect 396 395 397 396
tri 397 395 398 396 nw
tri 398 395 399 396 ne
rect 399 395 400 396
tri 400 395 403 398 sw
tri 390 392 393 395 se
tri 393 392 396 395 nw
tri 400 392 403 395 ne
tri 403 392 406 395 sw
tri 390 390 392 392 ne
tri 392 390 393 392 nw
tri 403 390 404 392 ne
tri 404 390 406 392 nw
rect 466 330 467 343
tri 467 330 471 334 se
tri 530 330 534 334 sw
rect 534 330 535 343
rect 466 329 535 330
rect 466 317 467 329
tri 467 325 471 329 ne
tri 530 325 534 329 nw
rect 534 317 535 329
rect 669 330 670 343
tri 670 330 674 334 se
tri 765 330 769 334 sw
rect 769 330 770 343
rect 669 329 770 330
rect 669 317 670 329
tri 670 325 674 329 ne
tri 765 325 769 329 nw
rect 769 317 770 329
rect 189 176 190 189
tri 190 176 194 180 se
tri 602 176 606 180 sw
rect 606 176 607 189
rect 189 175 377 176
rect 419 175 607 176
rect 189 163 190 175
tri 190 171 194 175 ne
tri 602 171 606 175 nw
rect 606 163 607 175
rect 362 136 363 149
tri 363 136 367 140 se
tri 429 136 433 140 sw
rect 433 136 434 149
rect 362 135 434 136
rect 362 123 363 135
tri 363 131 367 135 ne
tri 429 131 433 135 nw
rect 433 123 434 135
<< labels >>
flabel comment s 405 90 405 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 405 223 405 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 169 517 169 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 169 496 169 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 397 148 397 148 0 FreeSans 100 0 0 0 0.360
flabel comment s 398 783 398 783 0 FreeSans 100 0 0 0 3.720
flabel comment s 398 621 398 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 719 342 719 342 0 FreeSans 100 0 0 0 0.505
flabel comment s 638 545 638 545 0 FreeSans 100 0 0 0 0.310
flabel comment s 224 454 224 454 0 FreeSans 100 0 0 0 0.360
flabel comment s 500 342 500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s 398 177 398 177 0 FreeSans 100 0 0 0 2.090
flabel comment s 398 480 398 480 0 FreeSans 100 0 0 0 0.068
<< properties >>
string GDS_END 8229068
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 8221600
<< end >>
