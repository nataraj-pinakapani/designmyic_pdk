magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< dnwell >>
rect 795 16049 2256 22957
rect 23661 569 25900 1239
<< nwell >>
rect 2150 23053 2454 25429
rect 710 22751 2454 23053
rect 710 16255 1012 22751
rect 2150 16255 2454 22751
rect 710 15953 2454 16255
rect 2150 15591 2454 15953
rect -57 13363 26923 13785
rect -57 5423 365 13363
rect 779 6526 26099 12963
rect 26501 5423 26923 13363
rect -57 5121 26923 5423
rect 6177 1542 8670 2783
rect 14929 2283 18183 2777
rect 24267 2451 24801 2783
rect 15690 1542 18183 2283
rect 23581 1033 25980 1319
rect 23581 775 23867 1033
rect 25694 775 25980 1033
rect 23581 489 25980 775
<< pwell >>
rect 1072 22537 1850 22691
rect 1072 22347 1226 22537
rect 1696 22347 1850 22537
rect 1072 20963 1850 22347
rect 1072 16490 1226 20963
rect 1696 16490 1850 20963
rect 1072 16336 1850 16490
rect 491 13026 26420 13248
rect 491 5877 713 13026
rect 26198 5877 26420 13026
rect 491 5655 26420 5877
rect 24307 2863 24585 3055
rect 23927 835 25629 971
<< mvnmos >>
rect 1333 21721 1433 22321
rect 1489 21721 1589 22321
rect 1333 20989 1433 21589
rect 1489 20989 1589 21589
rect 24386 2889 24506 3029
rect 24114 861 24214 945
rect 24270 861 24370 945
rect 24426 861 24526 945
rect 24582 861 24682 945
rect 24874 861 24974 945
rect 25030 861 25130 945
rect 25186 861 25286 945
rect 25342 861 25442 945
<< mvpmos >>
rect 1732 9895 1832 10495
rect 1888 9895 1988 10495
rect 1289 9099 1389 9699
rect 1445 9099 1545 9699
rect 6552 2633 6752 2717
rect 24386 2517 24506 2717
rect 24562 2517 24682 2717
<< mvndiff >>
rect 1280 22243 1333 22321
rect 1280 22209 1288 22243
rect 1322 22209 1333 22243
rect 1280 22175 1333 22209
rect 1280 22141 1288 22175
rect 1322 22141 1333 22175
rect 1280 22107 1333 22141
rect 1280 22073 1288 22107
rect 1322 22073 1333 22107
rect 1280 22039 1333 22073
rect 1280 22005 1288 22039
rect 1322 22005 1333 22039
rect 1280 21971 1333 22005
rect 1280 21937 1288 21971
rect 1322 21937 1333 21971
rect 1280 21903 1333 21937
rect 1280 21869 1288 21903
rect 1322 21869 1333 21903
rect 1280 21835 1333 21869
rect 1280 21801 1288 21835
rect 1322 21801 1333 21835
rect 1280 21767 1333 21801
rect 1280 21733 1288 21767
rect 1322 21733 1333 21767
rect 1280 21721 1333 21733
rect 1433 22243 1489 22321
rect 1433 22209 1444 22243
rect 1478 22209 1489 22243
rect 1433 22175 1489 22209
rect 1433 22141 1444 22175
rect 1478 22141 1489 22175
rect 1433 22107 1489 22141
rect 1433 22073 1444 22107
rect 1478 22073 1489 22107
rect 1433 22039 1489 22073
rect 1433 22005 1444 22039
rect 1478 22005 1489 22039
rect 1433 21971 1489 22005
rect 1433 21937 1444 21971
rect 1478 21937 1489 21971
rect 1433 21903 1489 21937
rect 1433 21869 1444 21903
rect 1478 21869 1489 21903
rect 1433 21835 1489 21869
rect 1433 21801 1444 21835
rect 1478 21801 1489 21835
rect 1433 21767 1489 21801
rect 1433 21733 1444 21767
rect 1478 21733 1489 21767
rect 1433 21721 1489 21733
rect 1589 22243 1642 22321
rect 1589 22209 1600 22243
rect 1634 22209 1642 22243
rect 1589 22175 1642 22209
rect 1589 22141 1600 22175
rect 1634 22141 1642 22175
rect 1589 22107 1642 22141
rect 1589 22073 1600 22107
rect 1634 22073 1642 22107
rect 1589 22039 1642 22073
rect 1589 22005 1600 22039
rect 1634 22005 1642 22039
rect 1589 21971 1642 22005
rect 1589 21937 1600 21971
rect 1634 21937 1642 21971
rect 1589 21903 1642 21937
rect 1589 21869 1600 21903
rect 1634 21869 1642 21903
rect 1589 21835 1642 21869
rect 1589 21801 1600 21835
rect 1634 21801 1642 21835
rect 1589 21767 1642 21801
rect 1589 21733 1600 21767
rect 1634 21733 1642 21767
rect 1589 21721 1642 21733
rect 1280 21577 1333 21589
rect 1280 21543 1288 21577
rect 1322 21543 1333 21577
rect 1280 21509 1333 21543
rect 1280 21475 1288 21509
rect 1322 21475 1333 21509
rect 1280 21441 1333 21475
rect 1280 21407 1288 21441
rect 1322 21407 1333 21441
rect 1280 21373 1333 21407
rect 1280 21339 1288 21373
rect 1322 21339 1333 21373
rect 1280 21305 1333 21339
rect 1280 21271 1288 21305
rect 1322 21271 1333 21305
rect 1280 21237 1333 21271
rect 1280 21203 1288 21237
rect 1322 21203 1333 21237
rect 1280 21169 1333 21203
rect 1280 21135 1288 21169
rect 1322 21135 1333 21169
rect 1280 21101 1333 21135
rect 1280 21067 1288 21101
rect 1322 21067 1333 21101
rect 1280 20989 1333 21067
rect 1433 21577 1489 21589
rect 1433 21543 1444 21577
rect 1478 21543 1489 21577
rect 1433 21509 1489 21543
rect 1433 21475 1444 21509
rect 1478 21475 1489 21509
rect 1433 21441 1489 21475
rect 1433 21407 1444 21441
rect 1478 21407 1489 21441
rect 1433 21373 1489 21407
rect 1433 21339 1444 21373
rect 1478 21339 1489 21373
rect 1433 21305 1489 21339
rect 1433 21271 1444 21305
rect 1478 21271 1489 21305
rect 1433 21237 1489 21271
rect 1433 21203 1444 21237
rect 1478 21203 1489 21237
rect 1433 21169 1489 21203
rect 1433 21135 1444 21169
rect 1478 21135 1489 21169
rect 1433 21101 1489 21135
rect 1433 21067 1444 21101
rect 1478 21067 1489 21101
rect 1433 20989 1489 21067
rect 1589 21577 1642 21589
rect 1589 21543 1600 21577
rect 1634 21543 1642 21577
rect 1589 21509 1642 21543
rect 1589 21475 1600 21509
rect 1634 21475 1642 21509
rect 1589 21441 1642 21475
rect 1589 21407 1600 21441
rect 1634 21407 1642 21441
rect 1589 21373 1642 21407
rect 1589 21339 1600 21373
rect 1634 21339 1642 21373
rect 1589 21305 1642 21339
rect 1589 21271 1600 21305
rect 1634 21271 1642 21305
rect 1589 21237 1642 21271
rect 1589 21203 1600 21237
rect 1634 21203 1642 21237
rect 1589 21169 1642 21203
rect 1589 21135 1600 21169
rect 1634 21135 1642 21169
rect 1589 21101 1642 21135
rect 1589 21067 1600 21101
rect 1634 21067 1642 21101
rect 1589 20989 1642 21067
rect 24333 3017 24386 3029
rect 24333 2983 24341 3017
rect 24375 2983 24386 3017
rect 24333 2949 24386 2983
rect 24333 2915 24341 2949
rect 24375 2915 24386 2949
rect 24333 2889 24386 2915
rect 24506 3017 24559 3029
rect 24506 2983 24517 3017
rect 24551 2983 24559 3017
rect 24506 2949 24559 2983
rect 24506 2915 24517 2949
rect 24551 2915 24559 2949
rect 24506 2889 24559 2915
rect 24061 933 24114 945
rect 24061 899 24069 933
rect 24103 899 24114 933
rect 24061 861 24114 899
rect 24214 933 24270 945
rect 24214 899 24225 933
rect 24259 899 24270 933
rect 24214 861 24270 899
rect 24370 933 24426 945
rect 24370 899 24381 933
rect 24415 899 24426 933
rect 24370 861 24426 899
rect 24526 933 24582 945
rect 24526 899 24537 933
rect 24571 899 24582 933
rect 24526 861 24582 899
rect 24682 933 24735 945
rect 24682 899 24693 933
rect 24727 899 24735 933
rect 24682 861 24735 899
rect 24821 907 24874 945
rect 24821 873 24829 907
rect 24863 873 24874 907
rect 24821 861 24874 873
rect 24974 907 25030 945
rect 24974 873 24985 907
rect 25019 873 25030 907
rect 24974 861 25030 873
rect 25130 907 25186 945
rect 25130 873 25141 907
rect 25175 873 25186 907
rect 25130 861 25186 873
rect 25286 907 25342 945
rect 25286 873 25297 907
rect 25331 873 25342 907
rect 25286 861 25342 873
rect 25442 907 25495 945
rect 25442 873 25453 907
rect 25487 873 25495 907
rect 25442 861 25495 873
<< mvpdiff >>
rect 1679 10483 1732 10495
rect 1679 10449 1687 10483
rect 1721 10449 1732 10483
rect 1679 10415 1732 10449
rect 1679 10381 1687 10415
rect 1721 10381 1732 10415
rect 1679 10347 1732 10381
rect 1679 10313 1687 10347
rect 1721 10313 1732 10347
rect 1679 10279 1732 10313
rect 1679 10245 1687 10279
rect 1721 10245 1732 10279
rect 1679 10211 1732 10245
rect 1679 10177 1687 10211
rect 1721 10177 1732 10211
rect 1679 10143 1732 10177
rect 1679 10109 1687 10143
rect 1721 10109 1732 10143
rect 1679 10075 1732 10109
rect 1679 10041 1687 10075
rect 1721 10041 1732 10075
rect 1679 10007 1732 10041
rect 1679 9973 1687 10007
rect 1721 9973 1732 10007
rect 1679 9895 1732 9973
rect 1832 10483 1888 10495
rect 1832 10449 1843 10483
rect 1877 10449 1888 10483
rect 1832 10415 1888 10449
rect 1832 10381 1843 10415
rect 1877 10381 1888 10415
rect 1832 10347 1888 10381
rect 1832 10313 1843 10347
rect 1877 10313 1888 10347
rect 1832 10279 1888 10313
rect 1832 10245 1843 10279
rect 1877 10245 1888 10279
rect 1832 10211 1888 10245
rect 1832 10177 1843 10211
rect 1877 10177 1888 10211
rect 1832 10143 1888 10177
rect 1832 10109 1843 10143
rect 1877 10109 1888 10143
rect 1832 10075 1888 10109
rect 1832 10041 1843 10075
rect 1877 10041 1888 10075
rect 1832 10007 1888 10041
rect 1832 9973 1843 10007
rect 1877 9973 1888 10007
rect 1832 9895 1888 9973
rect 1988 10483 2041 10495
rect 1988 10449 1999 10483
rect 2033 10449 2041 10483
rect 1988 10415 2041 10449
rect 1988 10381 1999 10415
rect 2033 10381 2041 10415
rect 1988 10347 2041 10381
rect 1988 10313 1999 10347
rect 2033 10313 2041 10347
rect 1988 10279 2041 10313
rect 1988 10245 1999 10279
rect 2033 10245 2041 10279
rect 1988 10211 2041 10245
rect 1988 10177 1999 10211
rect 2033 10177 2041 10211
rect 1988 10143 2041 10177
rect 1988 10109 1999 10143
rect 2033 10109 2041 10143
rect 1988 10075 2041 10109
rect 1988 10041 1999 10075
rect 2033 10041 2041 10075
rect 1988 10007 2041 10041
rect 1988 9973 1999 10007
rect 2033 9973 2041 10007
rect 1988 9895 2041 9973
rect 1236 9687 1289 9699
rect 1236 9653 1244 9687
rect 1278 9653 1289 9687
rect 1236 9619 1289 9653
rect 1236 9585 1244 9619
rect 1278 9585 1289 9619
rect 1236 9551 1289 9585
rect 1236 9517 1244 9551
rect 1278 9517 1289 9551
rect 1236 9483 1289 9517
rect 1236 9449 1244 9483
rect 1278 9449 1289 9483
rect 1236 9415 1289 9449
rect 1236 9381 1244 9415
rect 1278 9381 1289 9415
rect 1236 9347 1289 9381
rect 1236 9313 1244 9347
rect 1278 9313 1289 9347
rect 1236 9279 1289 9313
rect 1236 9245 1244 9279
rect 1278 9245 1289 9279
rect 1236 9211 1289 9245
rect 1236 9177 1244 9211
rect 1278 9177 1289 9211
rect 1236 9099 1289 9177
rect 1389 9687 1445 9699
rect 1389 9653 1400 9687
rect 1434 9653 1445 9687
rect 1389 9619 1445 9653
rect 1389 9585 1400 9619
rect 1434 9585 1445 9619
rect 1389 9551 1445 9585
rect 1389 9517 1400 9551
rect 1434 9517 1445 9551
rect 1389 9483 1445 9517
rect 1389 9449 1400 9483
rect 1434 9449 1445 9483
rect 1389 9415 1445 9449
rect 1389 9381 1400 9415
rect 1434 9381 1445 9415
rect 1389 9347 1445 9381
rect 1389 9313 1400 9347
rect 1434 9313 1445 9347
rect 1389 9279 1445 9313
rect 1389 9245 1400 9279
rect 1434 9245 1445 9279
rect 1389 9211 1445 9245
rect 1389 9177 1400 9211
rect 1434 9177 1445 9211
rect 1389 9099 1445 9177
rect 1545 9687 1598 9699
rect 1545 9653 1556 9687
rect 1590 9653 1598 9687
rect 1545 9619 1598 9653
rect 1545 9585 1556 9619
rect 1590 9585 1598 9619
rect 1545 9551 1598 9585
rect 1545 9517 1556 9551
rect 1590 9517 1598 9551
rect 1545 9483 1598 9517
rect 1545 9449 1556 9483
rect 1590 9449 1598 9483
rect 1545 9415 1598 9449
rect 1545 9381 1556 9415
rect 1590 9381 1598 9415
rect 1545 9347 1598 9381
rect 1545 9313 1556 9347
rect 1590 9313 1598 9347
rect 1545 9279 1598 9313
rect 1545 9245 1556 9279
rect 1590 9245 1598 9279
rect 1545 9211 1598 9245
rect 1545 9177 1556 9211
rect 1590 9177 1598 9211
rect 1545 9099 1598 9177
rect 6499 2705 6552 2717
rect 6499 2671 6507 2705
rect 6541 2671 6552 2705
rect 6499 2633 6552 2671
rect 6752 2705 6805 2717
rect 6752 2671 6763 2705
rect 6797 2671 6805 2705
rect 6752 2633 6805 2671
rect 24333 2699 24386 2717
rect 24333 2665 24341 2699
rect 24375 2665 24386 2699
rect 24333 2631 24386 2665
rect 24333 2597 24341 2631
rect 24375 2597 24386 2631
rect 24333 2563 24386 2597
rect 24333 2529 24341 2563
rect 24375 2529 24386 2563
rect 24333 2517 24386 2529
rect 24506 2699 24562 2717
rect 24506 2665 24517 2699
rect 24551 2665 24562 2699
rect 24506 2631 24562 2665
rect 24506 2597 24517 2631
rect 24551 2597 24562 2631
rect 24506 2563 24562 2597
rect 24506 2529 24517 2563
rect 24551 2529 24562 2563
rect 24506 2517 24562 2529
rect 24682 2699 24735 2717
rect 24682 2665 24693 2699
rect 24727 2665 24735 2699
rect 24682 2631 24735 2665
rect 24682 2597 24693 2631
rect 24727 2597 24735 2631
rect 24682 2563 24735 2597
rect 24682 2529 24693 2563
rect 24727 2529 24735 2563
rect 24682 2517 24735 2529
<< mvndiffc >>
rect 1288 22209 1322 22243
rect 1288 22141 1322 22175
rect 1288 22073 1322 22107
rect 1288 22005 1322 22039
rect 1288 21937 1322 21971
rect 1288 21869 1322 21903
rect 1288 21801 1322 21835
rect 1288 21733 1322 21767
rect 1444 22209 1478 22243
rect 1444 22141 1478 22175
rect 1444 22073 1478 22107
rect 1444 22005 1478 22039
rect 1444 21937 1478 21971
rect 1444 21869 1478 21903
rect 1444 21801 1478 21835
rect 1444 21733 1478 21767
rect 1600 22209 1634 22243
rect 1600 22141 1634 22175
rect 1600 22073 1634 22107
rect 1600 22005 1634 22039
rect 1600 21937 1634 21971
rect 1600 21869 1634 21903
rect 1600 21801 1634 21835
rect 1600 21733 1634 21767
rect 1288 21543 1322 21577
rect 1288 21475 1322 21509
rect 1288 21407 1322 21441
rect 1288 21339 1322 21373
rect 1288 21271 1322 21305
rect 1288 21203 1322 21237
rect 1288 21135 1322 21169
rect 1288 21067 1322 21101
rect 1444 21543 1478 21577
rect 1444 21475 1478 21509
rect 1444 21407 1478 21441
rect 1444 21339 1478 21373
rect 1444 21271 1478 21305
rect 1444 21203 1478 21237
rect 1444 21135 1478 21169
rect 1444 21067 1478 21101
rect 1600 21543 1634 21577
rect 1600 21475 1634 21509
rect 1600 21407 1634 21441
rect 1600 21339 1634 21373
rect 1600 21271 1634 21305
rect 1600 21203 1634 21237
rect 1600 21135 1634 21169
rect 1600 21067 1634 21101
rect 24341 2983 24375 3017
rect 24341 2915 24375 2949
rect 24517 2983 24551 3017
rect 24517 2915 24551 2949
rect 24069 899 24103 933
rect 24225 899 24259 933
rect 24381 899 24415 933
rect 24537 899 24571 933
rect 24693 899 24727 933
rect 24829 873 24863 907
rect 24985 873 25019 907
rect 25141 873 25175 907
rect 25297 873 25331 907
rect 25453 873 25487 907
<< mvpdiffc >>
rect 1687 10449 1721 10483
rect 1687 10381 1721 10415
rect 1687 10313 1721 10347
rect 1687 10245 1721 10279
rect 1687 10177 1721 10211
rect 1687 10109 1721 10143
rect 1687 10041 1721 10075
rect 1687 9973 1721 10007
rect 1843 10449 1877 10483
rect 1843 10381 1877 10415
rect 1843 10313 1877 10347
rect 1843 10245 1877 10279
rect 1843 10177 1877 10211
rect 1843 10109 1877 10143
rect 1843 10041 1877 10075
rect 1843 9973 1877 10007
rect 1999 10449 2033 10483
rect 1999 10381 2033 10415
rect 1999 10313 2033 10347
rect 1999 10245 2033 10279
rect 1999 10177 2033 10211
rect 1999 10109 2033 10143
rect 1999 10041 2033 10075
rect 1999 9973 2033 10007
rect 1244 9653 1278 9687
rect 1244 9585 1278 9619
rect 1244 9517 1278 9551
rect 1244 9449 1278 9483
rect 1244 9381 1278 9415
rect 1244 9313 1278 9347
rect 1244 9245 1278 9279
rect 1244 9177 1278 9211
rect 1400 9653 1434 9687
rect 1400 9585 1434 9619
rect 1400 9517 1434 9551
rect 1400 9449 1434 9483
rect 1400 9381 1434 9415
rect 1400 9313 1434 9347
rect 1400 9245 1434 9279
rect 1400 9177 1434 9211
rect 1556 9653 1590 9687
rect 1556 9585 1590 9619
rect 1556 9517 1590 9551
rect 1556 9449 1590 9483
rect 1556 9381 1590 9415
rect 1556 9313 1590 9347
rect 1556 9245 1590 9279
rect 1556 9177 1590 9211
rect 6507 2671 6541 2705
rect 6763 2671 6797 2705
rect 24341 2665 24375 2699
rect 24341 2597 24375 2631
rect 24341 2529 24375 2563
rect 24517 2665 24551 2699
rect 24517 2597 24551 2631
rect 24517 2529 24551 2563
rect 24693 2665 24727 2699
rect 24693 2597 24727 2631
rect 24693 2529 24727 2563
<< psubdiff >>
rect 1098 16749 1200 16778
rect 1098 16477 1200 16511
rect 1132 16464 1200 16477
rect 1132 16443 1166 16464
rect 1098 16362 1166 16443
rect 1676 16430 1722 16464
rect 1676 16396 1824 16430
rect 1676 16362 1710 16396
rect 1744 16362 1824 16396
<< mvpsubdiff >>
rect 1098 22631 1174 22665
rect 1208 22631 1314 22665
rect 1098 22597 1314 22631
rect 1200 22563 1314 22597
rect 1756 22584 1824 22665
rect 1756 22563 1790 22584
rect 1722 22550 1790 22563
rect 1722 22516 1824 22550
rect 1098 16778 1200 16783
rect 517 13154 585 13222
rect 551 13120 585 13154
rect 26119 13188 26154 13222
rect 26188 13188 26223 13222
rect 26257 13188 26292 13222
rect 26326 13188 26394 13222
rect 26119 13154 26394 13188
rect 26119 13120 26154 13154
rect 26188 13120 26223 13154
rect 26257 13120 26292 13154
rect 517 13085 653 13120
rect 551 13051 585 13085
rect 619 13052 653 13085
rect 26051 13086 26292 13120
rect 26051 13052 26086 13086
rect 26120 13052 26155 13086
rect 26189 13052 26224 13086
rect 619 13051 687 13052
rect 517 13017 687 13051
rect 517 13016 653 13017
rect 551 12982 585 13016
rect 619 12983 653 13016
rect 619 12982 687 12983
rect 517 12948 687 12982
rect 517 12947 653 12948
rect 551 12913 585 12947
rect 619 12914 653 12947
rect 619 12913 687 12914
rect 517 12879 687 12913
rect 517 12878 653 12879
rect 551 12844 585 12878
rect 619 12845 653 12878
rect 619 12844 687 12845
rect 517 12810 687 12844
rect 517 12809 653 12810
rect 551 12775 585 12809
rect 619 12776 653 12809
rect 619 12775 687 12776
rect 517 12741 687 12775
rect 517 12740 653 12741
rect 551 12706 585 12740
rect 619 12707 653 12740
rect 619 12706 687 12707
rect 517 12672 687 12706
rect 517 12671 653 12672
rect 551 12637 585 12671
rect 619 12638 653 12671
rect 619 12637 687 12638
rect 517 12603 687 12637
rect 517 12602 653 12603
rect 551 12568 585 12602
rect 619 12569 653 12602
rect 619 12568 687 12569
rect 517 12534 687 12568
rect 517 12533 653 12534
rect 551 12499 585 12533
rect 619 12500 653 12533
rect 619 12499 687 12500
rect 517 12465 687 12499
rect 517 12464 653 12465
rect 551 12430 585 12464
rect 619 12431 653 12464
rect 619 12430 687 12431
rect 517 12396 687 12430
rect 517 12395 653 12396
rect 551 12361 585 12395
rect 619 12362 653 12395
rect 619 12361 687 12362
rect 517 12327 687 12361
rect 517 12326 653 12327
rect 551 12292 585 12326
rect 619 12293 653 12326
rect 619 12292 687 12293
rect 517 12258 687 12292
rect 517 12257 653 12258
rect 551 12223 585 12257
rect 619 12224 653 12257
rect 619 12223 687 12224
rect 517 12189 687 12223
rect 517 12188 653 12189
rect 551 12154 585 12188
rect 619 12155 653 12188
rect 619 12154 687 12155
rect 517 12120 687 12154
rect 517 12119 653 12120
rect 551 12085 585 12119
rect 619 12086 653 12119
rect 619 12085 687 12086
rect 517 12051 687 12085
rect 517 12050 653 12051
rect 551 12016 585 12050
rect 619 12017 653 12050
rect 619 12016 687 12017
rect 517 11982 687 12016
rect 517 11981 653 11982
rect 551 11947 585 11981
rect 619 11948 653 11981
rect 619 11947 687 11948
rect 517 11913 687 11947
rect 517 11912 653 11913
rect 551 11878 585 11912
rect 619 11879 653 11912
rect 619 11878 687 11879
rect 517 11844 687 11878
rect 517 11843 653 11844
rect 551 11809 585 11843
rect 619 11810 653 11843
rect 619 11809 687 11810
rect 517 11775 687 11809
rect 517 11774 653 11775
rect 551 11740 585 11774
rect 619 11741 653 11774
rect 619 11740 687 11741
rect 517 11706 687 11740
rect 517 11705 653 11706
rect 551 11671 585 11705
rect 619 11672 653 11705
rect 619 11671 687 11672
rect 517 11637 687 11671
rect 517 11636 653 11637
rect 551 11602 585 11636
rect 619 11603 653 11636
rect 619 11602 687 11603
rect 517 11568 687 11602
rect 517 11567 653 11568
rect 551 11533 585 11567
rect 619 11534 653 11567
rect 619 11533 687 11534
rect 517 11499 687 11533
rect 517 11498 653 11499
rect 551 11464 585 11498
rect 619 11465 653 11498
rect 619 11464 687 11465
rect 517 11430 687 11464
rect 517 11429 653 11430
rect 551 11395 585 11429
rect 619 11396 653 11429
rect 619 11395 687 11396
rect 517 11361 687 11395
rect 517 11360 653 11361
rect 551 11326 585 11360
rect 619 11327 653 11360
rect 619 11326 687 11327
rect 517 11292 687 11326
rect 517 11291 653 11292
rect 551 11257 585 11291
rect 619 11258 653 11291
rect 619 11257 687 11258
rect 517 11223 687 11257
rect 517 11222 653 11223
rect 551 11188 585 11222
rect 619 11189 653 11222
rect 619 11188 687 11189
rect 517 11154 687 11188
rect 517 11153 653 11154
rect 551 11119 585 11153
rect 619 11120 653 11153
rect 619 11119 687 11120
rect 517 11085 687 11119
rect 517 11084 653 11085
rect 551 11050 585 11084
rect 619 11051 653 11084
rect 619 11050 687 11051
rect 517 11016 687 11050
rect 517 11015 653 11016
rect 551 10981 585 11015
rect 619 10982 653 11015
rect 619 10981 687 10982
rect 517 10947 687 10981
rect 517 10946 653 10947
rect 551 10912 585 10946
rect 619 10913 653 10946
rect 619 10912 687 10913
rect 517 10878 687 10912
rect 517 10877 653 10878
rect 551 10843 585 10877
rect 619 10844 653 10877
rect 619 10843 687 10844
rect 517 10809 687 10843
rect 517 10808 653 10809
rect 551 10774 585 10808
rect 619 10775 653 10808
rect 619 10774 687 10775
rect 517 10740 687 10774
rect 517 10739 653 10740
rect 551 10705 585 10739
rect 619 10706 653 10739
rect 619 10705 687 10706
rect 517 10671 687 10705
rect 517 10670 653 10671
rect 551 10636 585 10670
rect 619 10637 653 10670
rect 619 10636 687 10637
rect 517 10602 687 10636
rect 517 10601 653 10602
rect 551 10567 585 10601
rect 619 10568 653 10601
rect 619 10567 687 10568
rect 517 10533 687 10567
rect 517 10532 653 10533
rect 551 10498 585 10532
rect 619 10499 653 10532
rect 619 10498 687 10499
rect 517 10464 687 10498
rect 517 10463 653 10464
rect 551 10429 585 10463
rect 619 10430 653 10463
rect 619 10429 687 10430
rect 517 10395 687 10429
rect 517 10394 653 10395
rect 619 10361 653 10394
rect 619 10326 687 10361
rect 517 9748 687 9816
rect 551 9714 585 9748
rect 619 9714 653 9748
rect 517 9679 687 9714
rect 551 9645 585 9679
rect 619 9645 653 9679
rect 517 9610 687 9645
rect 551 9576 585 9610
rect 619 9576 653 9610
rect 517 9541 687 9576
rect 551 9507 585 9541
rect 619 9507 653 9541
rect 517 9472 687 9507
rect 551 9438 585 9472
rect 619 9438 653 9472
rect 517 9403 687 9438
rect 551 9369 585 9403
rect 619 9369 653 9403
rect 517 9334 687 9369
rect 551 9300 585 9334
rect 619 9300 653 9334
rect 517 9265 687 9300
rect 551 9231 585 9265
rect 619 9231 653 9265
rect 517 9196 687 9231
rect 551 9162 585 9196
rect 619 9162 653 9196
rect 517 9127 687 9162
rect 551 9093 585 9127
rect 619 9093 653 9127
rect 517 9058 687 9093
rect 551 9024 585 9058
rect 619 9024 653 9058
rect 517 8989 687 9024
rect 551 8955 585 8989
rect 619 8955 653 8989
rect 517 8920 687 8955
rect 551 8886 585 8920
rect 619 8886 653 8920
rect 517 8851 687 8886
rect 551 8817 585 8851
rect 619 8817 653 8851
rect 517 8782 687 8817
rect 551 8748 585 8782
rect 619 8748 653 8782
rect 517 8713 687 8748
rect 551 8679 585 8713
rect 619 8679 653 8713
rect 517 8644 687 8679
rect 551 8610 585 8644
rect 619 8610 653 8644
rect 517 8575 687 8610
rect 551 8541 585 8575
rect 619 8541 653 8575
rect 517 8506 687 8541
rect 551 8472 585 8506
rect 619 8472 653 8506
rect 517 8437 687 8472
rect 551 8403 585 8437
rect 619 8403 653 8437
rect 517 8368 687 8403
rect 551 8334 585 8368
rect 619 8334 653 8368
rect 517 8299 687 8334
rect 26224 7645 26292 7680
rect 26258 7612 26292 7645
rect 26258 7611 26394 7612
rect 26224 7577 26394 7611
rect 26224 7576 26292 7577
rect 26258 7543 26292 7576
rect 26326 7543 26360 7577
rect 26258 7542 26394 7543
rect 26224 7508 26394 7542
rect 26224 7507 26292 7508
rect 26258 7474 26292 7507
rect 26326 7474 26360 7508
rect 26258 7473 26394 7474
rect 26224 7439 26394 7473
rect 26224 7438 26292 7439
rect 26258 7405 26292 7438
rect 26326 7405 26360 7439
rect 26258 7404 26394 7405
rect 26224 7370 26394 7404
rect 26224 7369 26292 7370
rect 26258 7336 26292 7369
rect 26326 7336 26360 7370
rect 26258 7335 26394 7336
rect 26224 7301 26394 7335
rect 26224 7300 26292 7301
rect 26258 7267 26292 7300
rect 26326 7267 26360 7301
rect 26258 7266 26394 7267
rect 26224 7232 26394 7266
rect 26224 7231 26292 7232
rect 26258 7198 26292 7231
rect 26326 7198 26360 7232
rect 26258 7197 26394 7198
rect 26224 7163 26394 7197
rect 26224 7162 26292 7163
rect 26258 7129 26292 7162
rect 26326 7129 26360 7163
rect 26258 7128 26394 7129
rect 26224 7094 26394 7128
rect 26224 7093 26292 7094
rect 26258 7060 26292 7093
rect 26326 7060 26360 7094
rect 26258 7059 26394 7060
rect 26224 7025 26394 7059
rect 26224 7024 26292 7025
rect 26258 6991 26292 7024
rect 26326 6991 26360 7025
rect 26258 6990 26394 6991
rect 26224 6956 26394 6990
rect 26224 6955 26292 6956
rect 26258 6922 26292 6955
rect 26326 6922 26360 6956
rect 26258 6921 26394 6922
rect 26224 6887 26394 6921
rect 26224 6886 26292 6887
rect 26258 6853 26292 6886
rect 26326 6853 26360 6887
rect 26258 6852 26394 6853
rect 26224 6818 26394 6852
rect 26224 6817 26292 6818
rect 26258 6784 26292 6817
rect 26326 6784 26360 6818
rect 26258 6783 26394 6784
rect 26224 6749 26394 6783
rect 26224 6748 26292 6749
rect 26258 6715 26292 6748
rect 26326 6715 26360 6749
rect 26258 6714 26394 6715
rect 26224 6680 26394 6714
rect 26224 6679 26292 6680
rect 26258 6646 26292 6679
rect 26326 6646 26360 6680
rect 26258 6645 26394 6646
rect 26224 6611 26394 6645
rect 26224 6610 26292 6611
rect 26258 6577 26292 6610
rect 26326 6577 26360 6611
rect 26258 6576 26394 6577
rect 26224 6542 26394 6576
rect 26224 6541 26292 6542
rect 26258 6508 26292 6541
rect 26326 6508 26360 6542
rect 26258 6507 26394 6508
rect 26224 6473 26394 6507
rect 26224 6472 26292 6473
rect 26258 6439 26292 6472
rect 26326 6439 26360 6473
rect 26258 6438 26394 6439
rect 26224 6404 26394 6438
rect 26224 6403 26292 6404
rect 26258 6370 26292 6403
rect 26326 6370 26360 6404
rect 26258 6369 26394 6370
rect 26224 6335 26394 6369
rect 26224 6334 26292 6335
rect 26258 6301 26292 6334
rect 26326 6301 26360 6335
rect 26258 6300 26394 6301
rect 26224 6266 26394 6300
rect 26224 6265 26292 6266
rect 26258 6232 26292 6265
rect 26326 6232 26360 6266
rect 26258 6231 26394 6232
rect 26224 6197 26394 6231
rect 26224 6196 26292 6197
rect 26258 6163 26292 6196
rect 26326 6163 26360 6197
rect 26258 6162 26394 6163
rect 26224 6128 26394 6162
rect 26224 6127 26292 6128
rect 26258 6094 26292 6127
rect 26326 6094 26360 6128
rect 26258 6093 26394 6094
rect 26224 6059 26394 6093
rect 26224 6058 26292 6059
rect 26258 6025 26292 6058
rect 26326 6025 26360 6059
rect 26258 6024 26394 6025
rect 26224 5990 26394 6024
rect 26224 5989 26292 5990
rect 26258 5956 26292 5989
rect 26326 5956 26360 5990
rect 26258 5955 26394 5956
rect 26224 5921 26394 5955
rect 26224 5920 26292 5921
rect 26258 5887 26292 5920
rect 26326 5887 26360 5921
rect 26258 5886 26394 5887
rect 26224 5852 26394 5886
rect 26224 5851 26292 5852
rect 687 5817 722 5851
rect 756 5817 791 5851
rect 825 5817 860 5851
rect 619 5783 860 5817
rect 26258 5818 26292 5851
rect 26326 5818 26360 5852
rect 26258 5783 26394 5818
rect 619 5749 654 5783
rect 688 5749 723 5783
rect 757 5749 792 5783
rect 517 5715 792 5749
rect 517 5681 585 5715
rect 619 5681 654 5715
rect 688 5681 723 5715
rect 757 5681 792 5715
rect 26326 5749 26360 5783
rect 26326 5681 26394 5749
rect 23953 919 23987 945
rect 23953 861 23987 885
rect 25569 919 25603 945
rect 25569 861 25603 885
<< mvnsubdiff >>
rect 2217 25395 2387 25429
rect 776 22919 844 22987
rect 810 22885 844 22919
rect 1286 22953 1321 22987
rect 1355 22953 1390 22987
rect 1424 22953 1459 22987
rect 1493 22953 1528 22987
rect 1562 22953 1597 22987
rect 1631 22953 1666 22987
rect 1700 22953 1735 22987
rect 1769 22953 1804 22987
rect 1838 22953 1873 22987
rect 1907 22953 1942 22987
rect 1976 22953 2011 22987
rect 2045 22953 2080 22987
rect 2114 22953 2149 22987
rect 1286 22919 2149 22953
rect 1286 22885 1321 22919
rect 1355 22885 1390 22919
rect 1424 22885 1459 22919
rect 1493 22885 1528 22919
rect 1562 22885 1597 22919
rect 1631 22885 1666 22919
rect 1700 22885 1735 22919
rect 1769 22885 1804 22919
rect 1838 22885 1873 22919
rect 1907 22885 1942 22919
rect 1976 22885 2011 22919
rect 2045 22885 2080 22919
rect 2114 22885 2149 22919
rect 776 22850 912 22885
rect 810 22816 844 22850
rect 878 22817 912 22850
rect 1286 22851 2149 22885
rect 1286 22817 1321 22851
rect 1355 22817 1390 22851
rect 1424 22817 1459 22851
rect 1493 22817 1528 22851
rect 1562 22817 1597 22851
rect 1631 22817 1666 22851
rect 1700 22817 1735 22851
rect 1769 22817 1804 22851
rect 1838 22817 1873 22851
rect 1907 22817 1942 22851
rect 1976 22817 2011 22851
rect 2045 22817 2080 22851
rect 2114 22817 2149 22851
rect 878 22816 946 22817
rect 776 22782 946 22816
rect 776 22781 912 22782
rect 810 22747 844 22781
rect 878 22748 912 22781
rect 878 22747 946 22748
rect 776 22713 946 22747
rect 776 22712 912 22713
rect 810 22678 844 22712
rect 878 22679 912 22712
rect 878 22678 946 22679
rect 776 22644 946 22678
rect 776 22643 912 22644
rect 810 22609 844 22643
rect 878 22610 912 22643
rect 878 22609 946 22610
rect 776 22575 946 22609
rect 776 22574 912 22575
rect 810 22540 844 22574
rect 878 22541 912 22574
rect 878 22540 946 22541
rect 776 22506 946 22540
rect 776 22505 912 22506
rect 810 22471 844 22505
rect 878 22472 912 22505
rect 878 22471 946 22472
rect 776 22437 946 22471
rect 776 22436 912 22437
rect 810 22402 844 22436
rect 878 22403 912 22436
rect 878 22402 946 22403
rect 776 22368 946 22402
rect 776 22367 912 22368
rect 810 22333 844 22367
rect 878 22334 912 22367
rect 878 22333 946 22334
rect 776 22299 946 22333
rect 776 22298 912 22299
rect 810 22264 844 22298
rect 878 22265 912 22298
rect 878 22264 946 22265
rect 776 22230 946 22264
rect 776 22229 912 22230
rect 810 22195 844 22229
rect 878 22196 912 22229
rect 878 22195 946 22196
rect 776 22161 946 22195
rect 776 22160 912 22161
rect 810 22126 844 22160
rect 878 22127 912 22160
rect 878 22126 946 22127
rect 776 22092 946 22126
rect 776 22091 912 22092
rect 810 22057 844 22091
rect 878 22058 912 22091
rect 878 22057 946 22058
rect 776 22023 946 22057
rect 776 22022 912 22023
rect 810 21988 844 22022
rect 878 21989 912 22022
rect 878 21988 946 21989
rect 776 21954 946 21988
rect 776 21953 912 21954
rect 810 21919 844 21953
rect 878 21920 912 21953
rect 878 21919 946 21920
rect 776 21885 946 21919
rect 776 21884 912 21885
rect 810 21850 844 21884
rect 878 21851 912 21884
rect 878 21850 946 21851
rect 776 21816 946 21850
rect 776 21815 912 21816
rect 810 21781 844 21815
rect 878 21782 912 21815
rect 878 21781 946 21782
rect 776 21747 946 21781
rect 776 21746 912 21747
rect 810 21712 844 21746
rect 878 21713 912 21746
rect 878 21712 946 21713
rect 776 21678 946 21712
rect 776 21677 912 21678
rect 810 21643 844 21677
rect 878 21644 912 21677
rect 878 21643 946 21644
rect 776 21609 946 21643
rect 776 21608 912 21609
rect 810 21574 844 21608
rect 878 21575 912 21608
rect 878 21574 946 21575
rect 776 21540 946 21574
rect 776 21539 912 21540
rect 810 21505 844 21539
rect 878 21506 912 21539
rect 878 21505 946 21506
rect 776 21471 946 21505
rect 776 21470 912 21471
rect 810 21436 844 21470
rect 878 21437 912 21470
rect 878 21436 946 21437
rect 776 21402 946 21436
rect 776 21401 912 21402
rect 810 21367 844 21401
rect 878 21368 912 21401
rect 878 21367 946 21368
rect 776 21333 946 21367
rect 776 21332 912 21333
rect 810 21298 844 21332
rect 878 21299 912 21332
rect 878 21298 946 21299
rect 776 21264 946 21298
rect 776 21263 912 21264
rect 810 21229 844 21263
rect 878 21230 912 21263
rect 878 21229 946 21230
rect 776 21195 946 21229
rect 776 21194 912 21195
rect 810 21160 844 21194
rect 878 21161 912 21194
rect 878 21160 946 21161
rect 776 21126 946 21160
rect 776 21125 912 21126
rect 810 21091 844 21125
rect 878 21092 912 21125
rect 878 21091 946 21092
rect 776 21057 946 21091
rect 776 21056 912 21057
rect 810 21022 844 21056
rect 878 21023 912 21056
rect 878 21022 946 21023
rect 776 20988 946 21022
rect 776 20987 912 20988
rect 810 20953 844 20987
rect 878 20954 912 20987
rect 878 20953 946 20954
rect 776 20919 946 20953
rect 776 20918 912 20919
rect 810 20884 844 20918
rect 878 20885 912 20918
rect 878 20884 946 20885
rect 776 20850 946 20884
rect 776 20849 912 20850
rect 810 20815 844 20849
rect 878 20816 912 20849
rect 878 20815 946 20816
rect 776 20781 946 20815
rect 776 20780 912 20781
rect 810 20746 844 20780
rect 878 20747 912 20780
rect 878 20746 946 20747
rect 776 20712 946 20746
rect 776 20711 912 20712
rect 810 20677 844 20711
rect 878 20678 912 20711
rect 878 20677 946 20678
rect 776 20643 946 20677
rect 776 20642 912 20643
rect 810 20608 844 20642
rect 878 20609 912 20642
rect 878 20608 946 20609
rect 776 20574 946 20608
rect 776 20573 912 20574
rect 810 20539 844 20573
rect 878 20540 912 20573
rect 878 20539 946 20540
rect 776 20505 946 20539
rect 776 20504 912 20505
rect 810 20470 844 20504
rect 878 20471 912 20504
rect 878 20470 946 20471
rect 776 20436 946 20470
rect 776 20435 912 20436
rect 810 20401 844 20435
rect 878 20402 912 20435
rect 878 20401 946 20402
rect 776 20367 946 20401
rect 776 20366 912 20367
rect 810 20332 844 20366
rect 878 20333 912 20366
rect 878 20332 946 20333
rect 776 20298 946 20332
rect 776 20297 912 20298
rect 810 20263 844 20297
rect 878 20264 912 20297
rect 878 20263 946 20264
rect 776 20229 946 20263
rect 776 20228 912 20229
rect 810 20194 844 20228
rect 878 20195 912 20228
rect 878 20194 946 20195
rect 776 20160 946 20194
rect 776 20159 912 20160
rect 810 20125 844 20159
rect 878 20126 912 20159
rect 878 20125 946 20126
rect 776 20091 946 20125
rect 776 20090 912 20091
rect 810 20056 844 20090
rect 878 20057 912 20090
rect 878 20056 946 20057
rect 776 20022 946 20056
rect 776 20021 912 20022
rect 810 19987 844 20021
rect 878 19988 912 20021
rect 878 19987 946 19988
rect 776 19953 946 19987
rect 776 19952 912 19953
rect 810 19918 844 19952
rect 878 19919 912 19952
rect 878 19918 946 19919
rect 776 19884 946 19918
rect 776 19883 912 19884
rect 810 19849 844 19883
rect 878 19850 912 19883
rect 878 19849 946 19850
rect 776 19815 946 19849
rect 776 19814 912 19815
rect 810 19780 844 19814
rect 878 19781 912 19814
rect 878 19780 946 19781
rect 776 19746 946 19780
rect 776 19745 912 19746
rect 810 19711 844 19745
rect 878 19712 912 19745
rect 878 19711 946 19712
rect 776 19677 946 19711
rect 776 19676 912 19677
rect 810 19642 844 19676
rect 878 19643 912 19676
rect 878 19642 946 19643
rect 776 19608 946 19642
rect 776 19607 912 19608
rect 810 19573 844 19607
rect 878 19574 912 19607
rect 878 19573 946 19574
rect 776 19539 946 19573
rect 776 19538 912 19539
rect 810 19504 844 19538
rect 878 19505 912 19538
rect 878 19504 946 19505
rect 776 19470 946 19504
rect 776 19469 912 19470
rect 810 19435 844 19469
rect 878 19436 912 19469
rect 878 19435 946 19436
rect 776 19401 946 19435
rect 776 19400 912 19401
rect 810 19366 844 19400
rect 878 19367 912 19400
rect 878 19366 946 19367
rect 776 19332 946 19366
rect 776 19331 912 19332
rect 810 19297 844 19331
rect 878 19298 912 19331
rect 878 19297 946 19298
rect 776 19263 946 19297
rect 776 19262 912 19263
rect 810 19228 844 19262
rect 878 19229 912 19262
rect 878 19228 946 19229
rect 776 19194 946 19228
rect 776 19193 912 19194
rect 810 19159 844 19193
rect 878 19160 912 19193
rect 878 19159 946 19160
rect 776 19125 946 19159
rect 776 19124 912 19125
rect 810 19090 844 19124
rect 878 19091 912 19124
rect 878 19090 946 19091
rect 776 19056 946 19090
rect 776 19055 912 19056
rect 810 19021 844 19055
rect 878 19022 912 19055
rect 878 19021 946 19022
rect 776 18987 946 19021
rect 776 18986 912 18987
rect 810 18952 844 18986
rect 878 18953 912 18986
rect 878 18952 946 18953
rect 776 18918 946 18952
rect 776 18917 912 18918
rect 810 18883 844 18917
rect 878 18884 912 18917
rect 878 18883 946 18884
rect 776 18849 946 18883
rect 776 18848 912 18849
rect 810 18814 844 18848
rect 878 18815 912 18848
rect 878 18814 946 18815
rect 776 18780 946 18814
rect 776 18779 912 18780
rect 810 18745 844 18779
rect 878 18746 912 18779
rect 878 18745 946 18746
rect 776 18711 946 18745
rect 776 18710 912 18711
rect 810 18676 844 18710
rect 878 18677 912 18710
rect 878 18676 946 18677
rect 776 18642 946 18676
rect 776 18641 912 18642
rect 810 18607 844 18641
rect 878 18608 912 18641
rect 878 18607 946 18608
rect 776 18573 946 18607
rect 776 18572 912 18573
rect 810 18538 844 18572
rect 878 18539 912 18572
rect 878 18538 946 18539
rect 776 18504 946 18538
rect 776 18503 912 18504
rect 810 18469 844 18503
rect 878 18470 912 18503
rect 878 18469 946 18470
rect 776 18435 946 18469
rect 776 18434 912 18435
rect 810 18400 844 18434
rect 878 18401 912 18434
rect 878 18400 946 18401
rect 776 18366 946 18400
rect 776 18365 912 18366
rect 878 18332 912 18365
rect 878 18297 946 18332
rect 2217 16418 2387 16453
rect 2251 16384 2285 16418
rect 2319 16384 2353 16418
rect 2217 16349 2387 16384
rect 2251 16315 2285 16349
rect 2319 16315 2353 16349
rect 2217 16280 2387 16315
rect 2251 16246 2285 16280
rect 2319 16246 2353 16280
rect 2217 16211 2387 16246
rect 946 16155 981 16189
rect 1015 16155 1050 16189
rect 1084 16155 1119 16189
rect 1153 16155 1188 16189
rect 1222 16155 1257 16189
rect 1291 16155 1326 16189
rect 1360 16155 1395 16189
rect 1429 16155 1464 16189
rect 1498 16155 1533 16189
rect 1567 16155 1602 16189
rect 1636 16155 1671 16189
rect 1705 16155 1740 16189
rect 1774 16155 1809 16189
rect 878 16121 1809 16155
rect 2183 16177 2217 16189
rect 2251 16177 2285 16211
rect 2319 16177 2353 16211
rect 2183 16142 2387 16177
rect 878 16087 913 16121
rect 947 16087 982 16121
rect 1016 16087 1051 16121
rect 1085 16087 1120 16121
rect 1154 16087 1189 16121
rect 1223 16087 1258 16121
rect 1292 16087 1327 16121
rect 1361 16087 1396 16121
rect 1430 16087 1465 16121
rect 1499 16087 1534 16121
rect 1568 16087 1603 16121
rect 1637 16087 1672 16121
rect 1706 16087 1741 16121
rect 776 16053 1741 16087
rect 776 16019 844 16053
rect 878 16019 913 16053
rect 947 16019 982 16053
rect 1016 16019 1051 16053
rect 1085 16019 1120 16053
rect 1154 16019 1189 16053
rect 1223 16019 1258 16053
rect 1292 16019 1327 16053
rect 1361 16019 1396 16053
rect 1430 16019 1465 16053
rect 1499 16019 1534 16053
rect 1568 16019 1603 16053
rect 1637 16019 1672 16053
rect 1706 16019 1741 16053
rect 2183 16108 2217 16142
rect 2251 16108 2285 16142
rect 2319 16108 2353 16142
rect 2183 16073 2387 16108
rect 2183 16039 2217 16073
rect 2251 16039 2285 16073
rect 2319 16039 2353 16073
rect 2183 16019 2387 16039
rect 2217 16004 2387 16019
rect 2251 15970 2285 16004
rect 2319 15970 2353 16004
rect 2217 15935 2387 15970
rect 2251 15901 2285 15935
rect 2319 15901 2353 15935
rect 2217 15866 2387 15901
rect 2251 15832 2285 15866
rect 2319 15832 2353 15866
rect 2217 15797 2387 15832
rect 2251 15763 2285 15797
rect 2319 15763 2353 15797
rect 2217 15728 2387 15763
rect 2251 15694 2285 15728
rect 2319 15694 2353 15728
rect 2217 15659 2387 15694
rect 2251 15625 2285 15659
rect 2319 15625 2353 15659
rect 2217 15591 2387 15625
rect 69 13625 192 13659
rect 226 13625 260 13659
rect 69 13591 260 13625
rect 171 13557 260 13591
rect 171 13523 328 13557
rect 239 13489 328 13523
rect 26678 13489 26797 13659
rect 26627 13415 26797 13489
rect 903 12803 985 12837
rect 1019 12803 1053 12837
rect 903 12769 1053 12803
rect 1005 12735 1053 12769
rect 25907 12736 25975 12837
rect 25907 12735 25941 12736
rect 1005 12701 1121 12735
rect 1073 12667 1121 12701
rect 25839 12702 25941 12735
rect 25839 12668 25975 12702
rect 25839 12667 25873 12668
rect 25805 12600 25873 12667
rect 11355 8147 11505 8175
rect 11355 8113 11379 8147
rect 11413 8113 11447 8147
rect 11481 8113 11505 8147
rect 903 7169 1073 7295
rect 1005 6820 1073 6863
rect 1005 6795 1039 6820
rect 903 6761 1039 6795
rect 937 6752 1039 6761
rect 25757 6786 25805 6820
rect 25757 6752 25873 6786
rect 937 6727 971 6752
rect 903 6650 971 6727
rect 25825 6718 25873 6752
rect 25825 6684 25975 6718
rect 25825 6650 25859 6684
rect 25893 6650 25975 6684
rect 307 5323 342 5357
rect 376 5323 411 5357
rect 445 5323 480 5357
rect 514 5323 549 5357
rect 583 5323 618 5357
rect 652 5323 687 5357
rect 721 5323 756 5357
rect 790 5323 825 5357
rect 859 5323 894 5357
rect 928 5323 963 5357
rect 997 5323 1032 5357
rect 1066 5323 1101 5357
rect 1135 5323 1170 5357
rect 1204 5323 1239 5357
rect 1273 5323 1308 5357
rect 1342 5323 1377 5357
rect 1411 5323 1446 5357
rect 1480 5323 1515 5357
rect 1549 5323 1584 5357
rect 1618 5323 1653 5357
rect 1687 5323 1722 5357
rect 1756 5323 1791 5357
rect 1825 5323 1860 5357
rect 1894 5323 1929 5357
rect 1963 5323 1998 5357
rect 2032 5323 2067 5357
rect 2101 5323 2136 5357
rect 2170 5323 2205 5357
rect 2239 5323 2274 5357
rect 2308 5323 2343 5357
rect 2377 5323 2412 5357
rect 2446 5323 2481 5357
rect 2515 5323 2550 5357
rect 2584 5323 2619 5357
rect 2653 5323 2688 5357
rect 2722 5323 2757 5357
rect 2791 5323 2826 5357
rect 2860 5323 2895 5357
rect 307 5289 2895 5323
rect 69 5255 273 5261
rect 307 5255 342 5289
rect 376 5255 411 5289
rect 445 5255 480 5289
rect 514 5255 549 5289
rect 583 5255 618 5289
rect 652 5255 687 5289
rect 721 5255 756 5289
rect 790 5255 825 5289
rect 859 5255 894 5289
rect 928 5255 963 5289
rect 997 5255 1032 5289
rect 1066 5255 1101 5289
rect 1135 5255 1170 5289
rect 1204 5255 1239 5289
rect 1273 5255 1308 5289
rect 1342 5255 1377 5289
rect 1411 5255 1446 5289
rect 1480 5255 1515 5289
rect 1549 5255 1584 5289
rect 1618 5255 1653 5289
rect 1687 5255 1722 5289
rect 1756 5255 1791 5289
rect 1825 5255 1860 5289
rect 1894 5255 1929 5289
rect 1963 5255 1998 5289
rect 2032 5255 2067 5289
rect 2101 5255 2136 5289
rect 2170 5255 2205 5289
rect 2239 5255 2274 5289
rect 2308 5255 2343 5289
rect 2377 5255 2412 5289
rect 2446 5255 2481 5289
rect 2515 5255 2550 5289
rect 2584 5255 2619 5289
rect 2653 5255 2688 5289
rect 2722 5255 2757 5289
rect 2791 5255 2826 5289
rect 2860 5255 2895 5289
rect 69 5221 2895 5255
rect 69 5187 273 5221
rect 307 5187 342 5221
rect 376 5187 411 5221
rect 445 5187 480 5221
rect 514 5187 549 5221
rect 583 5187 618 5221
rect 652 5187 687 5221
rect 721 5187 756 5221
rect 790 5187 825 5221
rect 859 5187 894 5221
rect 928 5187 963 5221
rect 997 5187 1032 5221
rect 1066 5187 1101 5221
rect 1135 5187 1170 5221
rect 1204 5187 1239 5221
rect 1273 5187 1308 5221
rect 1342 5187 1377 5221
rect 1411 5187 1446 5221
rect 1480 5187 1515 5221
rect 1549 5187 1584 5221
rect 1618 5187 1653 5221
rect 1687 5187 1722 5221
rect 1756 5187 1791 5221
rect 1825 5187 1860 5221
rect 1894 5187 1929 5221
rect 1963 5187 1998 5221
rect 2032 5187 2067 5221
rect 2101 5187 2136 5221
rect 2170 5187 2205 5221
rect 2239 5187 2274 5221
rect 2308 5187 2343 5221
rect 2377 5187 2412 5221
rect 2446 5187 2481 5221
rect 2515 5187 2550 5221
rect 2584 5187 2619 5221
rect 2653 5187 2688 5221
rect 2722 5187 2757 5221
rect 2791 5187 2826 5221
rect 2860 5187 2895 5221
rect 26593 5187 26797 5221
rect 23707 1159 23780 1193
rect 23814 1159 23848 1193
rect 23882 1159 23916 1193
rect 23950 1159 23984 1193
rect 24018 1159 24052 1193
rect 24086 1159 24120 1193
rect 24154 1159 24188 1193
rect 24222 1159 24256 1193
rect 24290 1159 24324 1193
rect 24358 1159 24392 1193
rect 24426 1159 24460 1193
rect 24494 1159 24528 1193
rect 24562 1159 24596 1193
rect 24630 1159 24664 1193
rect 24698 1159 24732 1193
rect 24766 1159 24800 1193
rect 24834 1159 24868 1193
rect 24902 1159 24936 1193
rect 24970 1159 25004 1193
rect 25038 1159 25072 1193
rect 25106 1159 25140 1193
rect 25174 1159 25208 1193
rect 25242 1159 25276 1193
rect 25310 1159 25344 1193
rect 25378 1159 25412 1193
rect 25446 1159 25480 1193
rect 25514 1159 25548 1193
rect 25582 1159 25616 1193
rect 25650 1159 25684 1193
rect 25718 1159 25752 1193
rect 25786 1159 25854 1193
rect 23707 1125 23741 1159
rect 23707 1057 23741 1091
rect 25820 1125 25854 1159
rect 25820 1057 25854 1091
rect 23707 989 23741 1023
rect 23707 921 23741 955
rect 25820 989 25854 1023
rect 23707 853 23741 887
rect 25820 921 25854 955
rect 25820 853 25854 887
rect 23707 785 23741 819
rect 23707 649 23741 751
rect 25820 785 25854 819
rect 25820 717 25854 751
rect 25820 649 25854 683
rect 23707 615 23775 649
rect 23809 615 23843 649
rect 23877 615 23911 649
rect 23945 615 23979 649
rect 24013 615 24047 649
rect 24081 615 24115 649
rect 24149 615 24183 649
rect 24217 615 24251 649
rect 24285 615 24319 649
rect 24353 615 24387 649
rect 24421 615 24455 649
rect 24489 615 24523 649
rect 24557 615 24591 649
rect 24625 615 24659 649
rect 24693 615 24727 649
rect 24761 615 24795 649
rect 24829 615 24863 649
rect 24897 615 24931 649
rect 24965 615 24999 649
rect 25033 615 25067 649
rect 25101 615 25135 649
rect 25169 615 25203 649
rect 25237 615 25271 649
rect 25305 615 25339 649
rect 25373 615 25407 649
rect 25441 615 25475 649
rect 25509 615 25543 649
rect 25577 615 25611 649
rect 25645 615 25679 649
rect 25713 615 25747 649
rect 25781 615 25854 649
<< psubdiffcont >>
rect 1098 16511 1200 16749
rect 1098 16443 1132 16477
rect 1166 16362 1676 16464
rect 1722 16430 1824 16778
rect 1710 16362 1744 16396
<< mvpsubdiffcont >>
rect 1174 22631 1208 22665
rect 1098 16783 1200 22597
rect 1314 22563 1756 22665
rect 1790 22550 1824 22584
rect 1722 16778 1824 22516
rect 517 13120 551 13154
rect 585 13120 26119 13222
rect 26154 13188 26188 13222
rect 26223 13188 26257 13222
rect 26292 13188 26326 13222
rect 26154 13120 26188 13154
rect 26223 13120 26257 13154
rect 517 13051 551 13085
rect 585 13051 619 13085
rect 653 13052 26051 13120
rect 26292 13086 26394 13154
rect 26086 13052 26120 13086
rect 26155 13052 26189 13086
rect 517 12982 551 13016
rect 585 12982 619 13016
rect 653 12983 687 13017
rect 517 12913 551 12947
rect 585 12913 619 12947
rect 653 12914 687 12948
rect 517 12844 551 12878
rect 585 12844 619 12878
rect 653 12845 687 12879
rect 517 12775 551 12809
rect 585 12775 619 12809
rect 653 12776 687 12810
rect 517 12706 551 12740
rect 585 12706 619 12740
rect 653 12707 687 12741
rect 517 12637 551 12671
rect 585 12637 619 12671
rect 653 12638 687 12672
rect 517 12568 551 12602
rect 585 12568 619 12602
rect 653 12569 687 12603
rect 517 12499 551 12533
rect 585 12499 619 12533
rect 653 12500 687 12534
rect 517 12430 551 12464
rect 585 12430 619 12464
rect 653 12431 687 12465
rect 517 12361 551 12395
rect 585 12361 619 12395
rect 653 12362 687 12396
rect 517 12292 551 12326
rect 585 12292 619 12326
rect 653 12293 687 12327
rect 517 12223 551 12257
rect 585 12223 619 12257
rect 653 12224 687 12258
rect 517 12154 551 12188
rect 585 12154 619 12188
rect 653 12155 687 12189
rect 517 12085 551 12119
rect 585 12085 619 12119
rect 653 12086 687 12120
rect 517 12016 551 12050
rect 585 12016 619 12050
rect 653 12017 687 12051
rect 517 11947 551 11981
rect 585 11947 619 11981
rect 653 11948 687 11982
rect 517 11878 551 11912
rect 585 11878 619 11912
rect 653 11879 687 11913
rect 517 11809 551 11843
rect 585 11809 619 11843
rect 653 11810 687 11844
rect 517 11740 551 11774
rect 585 11740 619 11774
rect 653 11741 687 11775
rect 517 11671 551 11705
rect 585 11671 619 11705
rect 653 11672 687 11706
rect 517 11602 551 11636
rect 585 11602 619 11636
rect 653 11603 687 11637
rect 517 11533 551 11567
rect 585 11533 619 11567
rect 653 11534 687 11568
rect 517 11464 551 11498
rect 585 11464 619 11498
rect 653 11465 687 11499
rect 517 11395 551 11429
rect 585 11395 619 11429
rect 653 11396 687 11430
rect 517 11326 551 11360
rect 585 11326 619 11360
rect 653 11327 687 11361
rect 517 11257 551 11291
rect 585 11257 619 11291
rect 653 11258 687 11292
rect 517 11188 551 11222
rect 585 11188 619 11222
rect 653 11189 687 11223
rect 517 11119 551 11153
rect 585 11119 619 11153
rect 653 11120 687 11154
rect 517 11050 551 11084
rect 585 11050 619 11084
rect 653 11051 687 11085
rect 517 10981 551 11015
rect 585 10981 619 11015
rect 653 10982 687 11016
rect 517 10912 551 10946
rect 585 10912 619 10946
rect 653 10913 687 10947
rect 517 10843 551 10877
rect 585 10843 619 10877
rect 653 10844 687 10878
rect 517 10774 551 10808
rect 585 10774 619 10808
rect 653 10775 687 10809
rect 517 10705 551 10739
rect 585 10705 619 10739
rect 653 10706 687 10740
rect 517 10636 551 10670
rect 585 10636 619 10670
rect 653 10637 687 10671
rect 517 10567 551 10601
rect 585 10567 619 10601
rect 653 10568 687 10602
rect 517 10498 551 10532
rect 585 10498 619 10532
rect 653 10499 687 10533
rect 517 10429 551 10463
rect 585 10429 619 10463
rect 653 10430 687 10464
rect 517 10326 619 10394
rect 653 10361 687 10395
rect 517 9816 687 10326
rect 517 9714 551 9748
rect 585 9714 619 9748
rect 653 9714 687 9748
rect 517 9645 551 9679
rect 585 9645 619 9679
rect 653 9645 687 9679
rect 517 9576 551 9610
rect 585 9576 619 9610
rect 653 9576 687 9610
rect 517 9507 551 9541
rect 585 9507 619 9541
rect 653 9507 687 9541
rect 517 9438 551 9472
rect 585 9438 619 9472
rect 653 9438 687 9472
rect 517 9369 551 9403
rect 585 9369 619 9403
rect 653 9369 687 9403
rect 517 9300 551 9334
rect 585 9300 619 9334
rect 653 9300 687 9334
rect 517 9231 551 9265
rect 585 9231 619 9265
rect 653 9231 687 9265
rect 517 9162 551 9196
rect 585 9162 619 9196
rect 653 9162 687 9196
rect 517 9093 551 9127
rect 585 9093 619 9127
rect 653 9093 687 9127
rect 517 9024 551 9058
rect 585 9024 619 9058
rect 653 9024 687 9058
rect 517 8955 551 8989
rect 585 8955 619 8989
rect 653 8955 687 8989
rect 517 8886 551 8920
rect 585 8886 619 8920
rect 653 8886 687 8920
rect 517 8817 551 8851
rect 585 8817 619 8851
rect 653 8817 687 8851
rect 517 8748 551 8782
rect 585 8748 619 8782
rect 653 8748 687 8782
rect 517 8679 551 8713
rect 585 8679 619 8713
rect 653 8679 687 8713
rect 517 8610 551 8644
rect 585 8610 619 8644
rect 653 8610 687 8644
rect 517 8541 551 8575
rect 585 8541 619 8575
rect 653 8541 687 8575
rect 517 8472 551 8506
rect 585 8472 619 8506
rect 653 8472 687 8506
rect 517 8403 551 8437
rect 585 8403 619 8437
rect 653 8403 687 8437
rect 517 8334 551 8368
rect 585 8334 619 8368
rect 653 8334 687 8368
rect 517 5817 687 8299
rect 26224 7680 26394 13086
rect 26224 7611 26258 7645
rect 26292 7612 26394 7680
rect 26224 7542 26258 7576
rect 26292 7543 26326 7577
rect 26360 7543 26394 7577
rect 26224 7473 26258 7507
rect 26292 7474 26326 7508
rect 26360 7474 26394 7508
rect 26224 7404 26258 7438
rect 26292 7405 26326 7439
rect 26360 7405 26394 7439
rect 26224 7335 26258 7369
rect 26292 7336 26326 7370
rect 26360 7336 26394 7370
rect 26224 7266 26258 7300
rect 26292 7267 26326 7301
rect 26360 7267 26394 7301
rect 26224 7197 26258 7231
rect 26292 7198 26326 7232
rect 26360 7198 26394 7232
rect 26224 7128 26258 7162
rect 26292 7129 26326 7163
rect 26360 7129 26394 7163
rect 26224 7059 26258 7093
rect 26292 7060 26326 7094
rect 26360 7060 26394 7094
rect 26224 6990 26258 7024
rect 26292 6991 26326 7025
rect 26360 6991 26394 7025
rect 26224 6921 26258 6955
rect 26292 6922 26326 6956
rect 26360 6922 26394 6956
rect 26224 6852 26258 6886
rect 26292 6853 26326 6887
rect 26360 6853 26394 6887
rect 26224 6783 26258 6817
rect 26292 6784 26326 6818
rect 26360 6784 26394 6818
rect 26224 6714 26258 6748
rect 26292 6715 26326 6749
rect 26360 6715 26394 6749
rect 26224 6645 26258 6679
rect 26292 6646 26326 6680
rect 26360 6646 26394 6680
rect 26224 6576 26258 6610
rect 26292 6577 26326 6611
rect 26360 6577 26394 6611
rect 26224 6507 26258 6541
rect 26292 6508 26326 6542
rect 26360 6508 26394 6542
rect 26224 6438 26258 6472
rect 26292 6439 26326 6473
rect 26360 6439 26394 6473
rect 26224 6369 26258 6403
rect 26292 6370 26326 6404
rect 26360 6370 26394 6404
rect 26224 6300 26258 6334
rect 26292 6301 26326 6335
rect 26360 6301 26394 6335
rect 26224 6231 26258 6265
rect 26292 6232 26326 6266
rect 26360 6232 26394 6266
rect 26224 6162 26258 6196
rect 26292 6163 26326 6197
rect 26360 6163 26394 6197
rect 26224 6093 26258 6127
rect 26292 6094 26326 6128
rect 26360 6094 26394 6128
rect 26224 6024 26258 6058
rect 26292 6025 26326 6059
rect 26360 6025 26394 6059
rect 26224 5955 26258 5989
rect 26292 5956 26326 5990
rect 26360 5956 26394 5990
rect 26224 5886 26258 5920
rect 26292 5887 26326 5921
rect 26360 5887 26394 5921
rect 722 5817 756 5851
rect 791 5817 825 5851
rect 517 5749 619 5817
rect 860 5783 26258 5851
rect 26292 5818 26326 5852
rect 26360 5818 26394 5852
rect 654 5749 688 5783
rect 723 5749 757 5783
rect 585 5681 619 5715
rect 654 5681 688 5715
rect 723 5681 757 5715
rect 792 5681 26326 5783
rect 26360 5749 26394 5783
rect 23953 885 23987 919
rect 25569 885 25603 919
<< mvnsubdiffcont >>
rect 2217 22987 2387 25395
rect 776 22885 810 22919
rect 844 22885 1286 22987
rect 1321 22953 1355 22987
rect 1390 22953 1424 22987
rect 1459 22953 1493 22987
rect 1528 22953 1562 22987
rect 1597 22953 1631 22987
rect 1666 22953 1700 22987
rect 1735 22953 1769 22987
rect 1804 22953 1838 22987
rect 1873 22953 1907 22987
rect 1942 22953 1976 22987
rect 2011 22953 2045 22987
rect 2080 22953 2114 22987
rect 1321 22885 1355 22919
rect 1390 22885 1424 22919
rect 1459 22885 1493 22919
rect 1528 22885 1562 22919
rect 1597 22885 1631 22919
rect 1666 22885 1700 22919
rect 1735 22885 1769 22919
rect 1804 22885 1838 22919
rect 1873 22885 1907 22919
rect 1942 22885 1976 22919
rect 2011 22885 2045 22919
rect 2080 22885 2114 22919
rect 776 22816 810 22850
rect 844 22816 878 22850
rect 912 22817 1286 22885
rect 1321 22817 1355 22851
rect 1390 22817 1424 22851
rect 1459 22817 1493 22851
rect 1528 22817 1562 22851
rect 1597 22817 1631 22851
rect 1666 22817 1700 22851
rect 1735 22817 1769 22851
rect 1804 22817 1838 22851
rect 1873 22817 1907 22851
rect 1942 22817 1976 22851
rect 2011 22817 2045 22851
rect 2080 22817 2114 22851
rect 2149 22817 2387 22987
rect 776 22747 810 22781
rect 844 22747 878 22781
rect 912 22748 946 22782
rect 776 22678 810 22712
rect 844 22678 878 22712
rect 912 22679 946 22713
rect 776 22609 810 22643
rect 844 22609 878 22643
rect 912 22610 946 22644
rect 776 22540 810 22574
rect 844 22540 878 22574
rect 912 22541 946 22575
rect 776 22471 810 22505
rect 844 22471 878 22505
rect 912 22472 946 22506
rect 776 22402 810 22436
rect 844 22402 878 22436
rect 912 22403 946 22437
rect 776 22333 810 22367
rect 844 22333 878 22367
rect 912 22334 946 22368
rect 776 22264 810 22298
rect 844 22264 878 22298
rect 912 22265 946 22299
rect 776 22195 810 22229
rect 844 22195 878 22229
rect 912 22196 946 22230
rect 776 22126 810 22160
rect 844 22126 878 22160
rect 912 22127 946 22161
rect 776 22057 810 22091
rect 844 22057 878 22091
rect 912 22058 946 22092
rect 776 21988 810 22022
rect 844 21988 878 22022
rect 912 21989 946 22023
rect 776 21919 810 21953
rect 844 21919 878 21953
rect 912 21920 946 21954
rect 776 21850 810 21884
rect 844 21850 878 21884
rect 912 21851 946 21885
rect 776 21781 810 21815
rect 844 21781 878 21815
rect 912 21782 946 21816
rect 776 21712 810 21746
rect 844 21712 878 21746
rect 912 21713 946 21747
rect 776 21643 810 21677
rect 844 21643 878 21677
rect 912 21644 946 21678
rect 776 21574 810 21608
rect 844 21574 878 21608
rect 912 21575 946 21609
rect 776 21505 810 21539
rect 844 21505 878 21539
rect 912 21506 946 21540
rect 776 21436 810 21470
rect 844 21436 878 21470
rect 912 21437 946 21471
rect 776 21367 810 21401
rect 844 21367 878 21401
rect 912 21368 946 21402
rect 776 21298 810 21332
rect 844 21298 878 21332
rect 912 21299 946 21333
rect 776 21229 810 21263
rect 844 21229 878 21263
rect 912 21230 946 21264
rect 776 21160 810 21194
rect 844 21160 878 21194
rect 912 21161 946 21195
rect 776 21091 810 21125
rect 844 21091 878 21125
rect 912 21092 946 21126
rect 776 21022 810 21056
rect 844 21022 878 21056
rect 912 21023 946 21057
rect 776 20953 810 20987
rect 844 20953 878 20987
rect 912 20954 946 20988
rect 776 20884 810 20918
rect 844 20884 878 20918
rect 912 20885 946 20919
rect 776 20815 810 20849
rect 844 20815 878 20849
rect 912 20816 946 20850
rect 776 20746 810 20780
rect 844 20746 878 20780
rect 912 20747 946 20781
rect 776 20677 810 20711
rect 844 20677 878 20711
rect 912 20678 946 20712
rect 776 20608 810 20642
rect 844 20608 878 20642
rect 912 20609 946 20643
rect 776 20539 810 20573
rect 844 20539 878 20573
rect 912 20540 946 20574
rect 776 20470 810 20504
rect 844 20470 878 20504
rect 912 20471 946 20505
rect 776 20401 810 20435
rect 844 20401 878 20435
rect 912 20402 946 20436
rect 776 20332 810 20366
rect 844 20332 878 20366
rect 912 20333 946 20367
rect 776 20263 810 20297
rect 844 20263 878 20297
rect 912 20264 946 20298
rect 776 20194 810 20228
rect 844 20194 878 20228
rect 912 20195 946 20229
rect 776 20125 810 20159
rect 844 20125 878 20159
rect 912 20126 946 20160
rect 776 20056 810 20090
rect 844 20056 878 20090
rect 912 20057 946 20091
rect 776 19987 810 20021
rect 844 19987 878 20021
rect 912 19988 946 20022
rect 776 19918 810 19952
rect 844 19918 878 19952
rect 912 19919 946 19953
rect 776 19849 810 19883
rect 844 19849 878 19883
rect 912 19850 946 19884
rect 776 19780 810 19814
rect 844 19780 878 19814
rect 912 19781 946 19815
rect 776 19711 810 19745
rect 844 19711 878 19745
rect 912 19712 946 19746
rect 776 19642 810 19676
rect 844 19642 878 19676
rect 912 19643 946 19677
rect 776 19573 810 19607
rect 844 19573 878 19607
rect 912 19574 946 19608
rect 776 19504 810 19538
rect 844 19504 878 19538
rect 912 19505 946 19539
rect 776 19435 810 19469
rect 844 19435 878 19469
rect 912 19436 946 19470
rect 776 19366 810 19400
rect 844 19366 878 19400
rect 912 19367 946 19401
rect 776 19297 810 19331
rect 844 19297 878 19331
rect 912 19298 946 19332
rect 776 19228 810 19262
rect 844 19228 878 19262
rect 912 19229 946 19263
rect 776 19159 810 19193
rect 844 19159 878 19193
rect 912 19160 946 19194
rect 776 19090 810 19124
rect 844 19090 878 19124
rect 912 19091 946 19125
rect 776 19021 810 19055
rect 844 19021 878 19055
rect 912 19022 946 19056
rect 776 18952 810 18986
rect 844 18952 878 18986
rect 912 18953 946 18987
rect 776 18883 810 18917
rect 844 18883 878 18917
rect 912 18884 946 18918
rect 776 18814 810 18848
rect 844 18814 878 18848
rect 912 18815 946 18849
rect 776 18745 810 18779
rect 844 18745 878 18779
rect 912 18746 946 18780
rect 776 18676 810 18710
rect 844 18676 878 18710
rect 912 18677 946 18711
rect 776 18607 810 18641
rect 844 18607 878 18641
rect 912 18608 946 18642
rect 776 18538 810 18572
rect 844 18538 878 18572
rect 912 18539 946 18573
rect 776 18469 810 18503
rect 844 18469 878 18503
rect 912 18470 946 18504
rect 776 18400 810 18434
rect 844 18400 878 18434
rect 912 18401 946 18435
rect 776 18297 878 18365
rect 912 18332 946 18366
rect 776 16155 946 18297
rect 2217 16453 2387 22817
rect 2217 16384 2251 16418
rect 2285 16384 2319 16418
rect 2353 16384 2387 16418
rect 2217 16315 2251 16349
rect 2285 16315 2319 16349
rect 2353 16315 2387 16349
rect 2217 16246 2251 16280
rect 2285 16246 2319 16280
rect 2353 16246 2387 16280
rect 981 16155 1015 16189
rect 1050 16155 1084 16189
rect 1119 16155 1153 16189
rect 1188 16155 1222 16189
rect 1257 16155 1291 16189
rect 1326 16155 1360 16189
rect 1395 16155 1429 16189
rect 1464 16155 1498 16189
rect 1533 16155 1567 16189
rect 1602 16155 1636 16189
rect 1671 16155 1705 16189
rect 1740 16155 1774 16189
rect 776 16087 878 16155
rect 1809 16121 2183 16189
rect 2217 16177 2251 16211
rect 2285 16177 2319 16211
rect 2353 16177 2387 16211
rect 913 16087 947 16121
rect 982 16087 1016 16121
rect 1051 16087 1085 16121
rect 1120 16087 1154 16121
rect 1189 16087 1223 16121
rect 1258 16087 1292 16121
rect 1327 16087 1361 16121
rect 1396 16087 1430 16121
rect 1465 16087 1499 16121
rect 1534 16087 1568 16121
rect 1603 16087 1637 16121
rect 1672 16087 1706 16121
rect 844 16019 878 16053
rect 913 16019 947 16053
rect 982 16019 1016 16053
rect 1051 16019 1085 16053
rect 1120 16019 1154 16053
rect 1189 16019 1223 16053
rect 1258 16019 1292 16053
rect 1327 16019 1361 16053
rect 1396 16019 1430 16053
rect 1465 16019 1499 16053
rect 1534 16019 1568 16053
rect 1603 16019 1637 16053
rect 1672 16019 1706 16053
rect 1741 16019 2183 16121
rect 2217 16108 2251 16142
rect 2285 16108 2319 16142
rect 2353 16108 2387 16142
rect 2217 16039 2251 16073
rect 2285 16039 2319 16073
rect 2353 16039 2387 16073
rect 2217 15970 2251 16004
rect 2285 15970 2319 16004
rect 2353 15970 2387 16004
rect 2217 15901 2251 15935
rect 2285 15901 2319 15935
rect 2353 15901 2387 15935
rect 2217 15832 2251 15866
rect 2285 15832 2319 15866
rect 2353 15832 2387 15866
rect 2217 15763 2251 15797
rect 2285 15763 2319 15797
rect 2353 15763 2387 15797
rect 2217 15694 2251 15728
rect 2285 15694 2319 15728
rect 2353 15694 2387 15728
rect 2217 15625 2251 15659
rect 2285 15625 2319 15659
rect 2353 15625 2387 15659
rect 192 13625 226 13659
rect 69 13523 171 13591
rect 260 13557 26678 13659
rect 69 5357 239 13523
rect 328 13489 26678 13557
rect 985 12803 1019 12837
rect 903 12701 1005 12769
rect 1053 12735 25907 12837
rect 903 7295 1073 12701
rect 1121 12667 25839 12735
rect 25941 12702 25975 12736
rect 25873 12600 25975 12668
rect 11379 8113 11413 8147
rect 11447 8113 11481 8147
rect 903 6863 1073 7169
rect 903 6795 1005 6863
rect 903 6727 937 6761
rect 1039 6752 25757 6820
rect 25805 6786 25975 12600
rect 971 6650 25825 6752
rect 25873 6718 25975 6786
rect 25859 6650 25893 6684
rect 26627 5357 26797 13415
rect 69 5261 307 5357
rect 342 5323 376 5357
rect 411 5323 445 5357
rect 480 5323 514 5357
rect 549 5323 583 5357
rect 618 5323 652 5357
rect 687 5323 721 5357
rect 756 5323 790 5357
rect 825 5323 859 5357
rect 894 5323 928 5357
rect 963 5323 997 5357
rect 1032 5323 1066 5357
rect 1101 5323 1135 5357
rect 1170 5323 1204 5357
rect 1239 5323 1273 5357
rect 1308 5323 1342 5357
rect 1377 5323 1411 5357
rect 1446 5323 1480 5357
rect 1515 5323 1549 5357
rect 1584 5323 1618 5357
rect 1653 5323 1687 5357
rect 1722 5323 1756 5357
rect 1791 5323 1825 5357
rect 1860 5323 1894 5357
rect 1929 5323 1963 5357
rect 1998 5323 2032 5357
rect 2067 5323 2101 5357
rect 2136 5323 2170 5357
rect 2205 5323 2239 5357
rect 2274 5323 2308 5357
rect 2343 5323 2377 5357
rect 2412 5323 2446 5357
rect 2481 5323 2515 5357
rect 2550 5323 2584 5357
rect 2619 5323 2653 5357
rect 2688 5323 2722 5357
rect 2757 5323 2791 5357
rect 2826 5323 2860 5357
rect 273 5255 307 5261
rect 342 5255 376 5289
rect 411 5255 445 5289
rect 480 5255 514 5289
rect 549 5255 583 5289
rect 618 5255 652 5289
rect 687 5255 721 5289
rect 756 5255 790 5289
rect 825 5255 859 5289
rect 894 5255 928 5289
rect 963 5255 997 5289
rect 1032 5255 1066 5289
rect 1101 5255 1135 5289
rect 1170 5255 1204 5289
rect 1239 5255 1273 5289
rect 1308 5255 1342 5289
rect 1377 5255 1411 5289
rect 1446 5255 1480 5289
rect 1515 5255 1549 5289
rect 1584 5255 1618 5289
rect 1653 5255 1687 5289
rect 1722 5255 1756 5289
rect 1791 5255 1825 5289
rect 1860 5255 1894 5289
rect 1929 5255 1963 5289
rect 1998 5255 2032 5289
rect 2067 5255 2101 5289
rect 2136 5255 2170 5289
rect 2205 5255 2239 5289
rect 2274 5255 2308 5289
rect 2343 5255 2377 5289
rect 2412 5255 2446 5289
rect 2481 5255 2515 5289
rect 2550 5255 2584 5289
rect 2619 5255 2653 5289
rect 2688 5255 2722 5289
rect 2757 5255 2791 5289
rect 2826 5255 2860 5289
rect 2895 5221 26797 5357
rect 273 5187 307 5221
rect 342 5187 376 5221
rect 411 5187 445 5221
rect 480 5187 514 5221
rect 549 5187 583 5221
rect 618 5187 652 5221
rect 687 5187 721 5221
rect 756 5187 790 5221
rect 825 5187 859 5221
rect 894 5187 928 5221
rect 963 5187 997 5221
rect 1032 5187 1066 5221
rect 1101 5187 1135 5221
rect 1170 5187 1204 5221
rect 1239 5187 1273 5221
rect 1308 5187 1342 5221
rect 1377 5187 1411 5221
rect 1446 5187 1480 5221
rect 1515 5187 1549 5221
rect 1584 5187 1618 5221
rect 1653 5187 1687 5221
rect 1722 5187 1756 5221
rect 1791 5187 1825 5221
rect 1860 5187 1894 5221
rect 1929 5187 1963 5221
rect 1998 5187 2032 5221
rect 2067 5187 2101 5221
rect 2136 5187 2170 5221
rect 2205 5187 2239 5221
rect 2274 5187 2308 5221
rect 2343 5187 2377 5221
rect 2412 5187 2446 5221
rect 2481 5187 2515 5221
rect 2550 5187 2584 5221
rect 2619 5187 2653 5221
rect 2688 5187 2722 5221
rect 2757 5187 2791 5221
rect 2826 5187 2860 5221
rect 2895 5187 26593 5221
rect 23780 1159 23814 1193
rect 23848 1159 23882 1193
rect 23916 1159 23950 1193
rect 23984 1159 24018 1193
rect 24052 1159 24086 1193
rect 24120 1159 24154 1193
rect 24188 1159 24222 1193
rect 24256 1159 24290 1193
rect 24324 1159 24358 1193
rect 24392 1159 24426 1193
rect 24460 1159 24494 1193
rect 24528 1159 24562 1193
rect 24596 1159 24630 1193
rect 24664 1159 24698 1193
rect 24732 1159 24766 1193
rect 24800 1159 24834 1193
rect 24868 1159 24902 1193
rect 24936 1159 24970 1193
rect 25004 1159 25038 1193
rect 25072 1159 25106 1193
rect 25140 1159 25174 1193
rect 25208 1159 25242 1193
rect 25276 1159 25310 1193
rect 25344 1159 25378 1193
rect 25412 1159 25446 1193
rect 25480 1159 25514 1193
rect 25548 1159 25582 1193
rect 25616 1159 25650 1193
rect 25684 1159 25718 1193
rect 25752 1159 25786 1193
rect 23707 1091 23741 1125
rect 23707 1023 23741 1057
rect 25820 1091 25854 1125
rect 23707 955 23741 989
rect 25820 1023 25854 1057
rect 25820 955 25854 989
rect 23707 887 23741 921
rect 25820 887 25854 921
rect 23707 819 23741 853
rect 23707 751 23741 785
rect 25820 819 25854 853
rect 25820 751 25854 785
rect 25820 683 25854 717
rect 23775 615 23809 649
rect 23843 615 23877 649
rect 23911 615 23945 649
rect 23979 615 24013 649
rect 24047 615 24081 649
rect 24115 615 24149 649
rect 24183 615 24217 649
rect 24251 615 24285 649
rect 24319 615 24353 649
rect 24387 615 24421 649
rect 24455 615 24489 649
rect 24523 615 24557 649
rect 24591 615 24625 649
rect 24659 615 24693 649
rect 24727 615 24761 649
rect 24795 615 24829 649
rect 24863 615 24897 649
rect 24931 615 24965 649
rect 24999 615 25033 649
rect 25067 615 25101 649
rect 25135 615 25169 649
rect 25203 615 25237 649
rect 25271 615 25305 649
rect 25339 615 25373 649
rect 25407 615 25441 649
rect 25475 615 25509 649
rect 25543 615 25577 649
rect 25611 615 25645 649
rect 25679 615 25713 649
rect 25747 615 25781 649
<< poly >>
rect 1333 22404 1433 22427
rect 1333 22370 1366 22404
rect 1400 22370 1433 22404
rect 1333 22321 1433 22370
rect 1489 22404 1589 22427
rect 1489 22370 1522 22404
rect 1556 22370 1589 22404
rect 1489 22321 1589 22370
rect 1333 21672 1433 21721
rect 1333 21638 1366 21672
rect 1400 21638 1433 21672
rect 1333 21589 1433 21638
rect 1489 21672 1589 21721
rect 1489 21638 1522 21672
rect 1556 21638 1589 21672
rect 1489 21589 1589 21638
rect 1333 20963 1433 20989
rect 1489 20963 1589 20989
rect 1732 10584 1988 10607
rect 1732 10550 1748 10584
rect 1782 10550 1843 10584
rect 1877 10550 1938 10584
rect 1972 10550 1988 10584
rect 1732 10527 1988 10550
rect 1732 10495 1832 10527
rect 1888 10495 1988 10527
rect 1732 9863 1832 9895
rect 1888 9863 1988 9895
rect 1289 9788 1545 9811
rect 1289 9754 1305 9788
rect 1339 9754 1400 9788
rect 1434 9754 1495 9788
rect 1529 9754 1545 9788
rect 1289 9731 1545 9754
rect 1289 9699 1389 9731
rect 1445 9699 1545 9731
rect 1289 9067 1389 9099
rect 1445 9067 1545 9099
rect 24386 3029 24506 3061
rect 24386 2857 24506 2889
rect 24386 2825 24682 2857
rect 24386 2791 24406 2825
rect 24440 2791 24480 2825
rect 24514 2791 24554 2825
rect 24588 2791 24628 2825
rect 24662 2791 24682 2825
rect 24386 2760 24682 2791
rect 6552 2717 6752 2743
rect 24386 2717 24506 2760
rect 24562 2717 24682 2760
rect 6552 2607 6752 2633
rect 24386 2491 24506 2517
rect 24562 2491 24682 2517
rect -1142 2188 -742 2204
rect -645 2188 -245 2204
rect -149 2188 251 2204
rect 347 2188 747 2204
rect 24114 1027 24370 1043
rect 24114 993 24130 1027
rect 24164 993 24225 1027
rect 24259 993 24320 1027
rect 24354 993 24370 1027
rect 24114 977 24370 993
rect 24114 945 24214 977
rect 24270 945 24370 977
rect 24426 1027 24682 1043
rect 24426 993 24442 1027
rect 24476 993 24537 1027
rect 24571 993 24632 1027
rect 24666 993 24682 1027
rect 24426 977 24682 993
rect 24426 945 24526 977
rect 24582 945 24682 977
rect 24874 1027 25130 1043
rect 24874 993 24890 1027
rect 24924 993 24985 1027
rect 25019 993 25080 1027
rect 25114 993 25130 1027
rect 24874 977 25130 993
rect 24874 945 24974 977
rect 25030 945 25130 977
rect 25186 1027 25442 1043
rect 25186 993 25202 1027
rect 25236 993 25297 1027
rect 25331 993 25392 1027
rect 25426 993 25442 1027
rect 25186 977 25442 993
rect 25186 945 25286 977
rect 25342 945 25442 977
rect 24114 829 24214 861
rect 24270 829 24370 861
rect 24426 829 24526 861
rect 24582 829 24682 861
rect 24874 829 24974 861
rect 25030 829 25130 861
rect 25186 829 25286 861
rect 25342 829 25442 861
<< polycont >>
rect 1366 22370 1400 22404
rect 1522 22370 1556 22404
rect 1366 21638 1400 21672
rect 1522 21638 1556 21672
rect 1748 10550 1782 10584
rect 1843 10550 1877 10584
rect 1938 10550 1972 10584
rect 1305 9754 1339 9788
rect 1400 9754 1434 9788
rect 1495 9754 1529 9788
rect 24406 2791 24440 2825
rect 24480 2791 24514 2825
rect 24554 2791 24588 2825
rect 24628 2791 24662 2825
rect 24130 993 24164 1027
rect 24225 993 24259 1027
rect 24320 993 24354 1027
rect 24442 993 24476 1027
rect 24537 993 24571 1027
rect 24632 993 24666 1027
rect 24890 993 24924 1027
rect 24985 993 25019 1027
rect 25080 993 25114 1027
rect 25202 993 25236 1027
rect 25297 993 25331 1027
rect 25392 993 25426 1027
<< locali >>
rect 2217 25395 2387 25429
rect 776 22919 844 22987
rect 810 22885 844 22919
rect 1286 22953 1321 22987
rect 1355 22953 1390 22987
rect 1424 22953 1459 22987
rect 1493 22953 1528 22987
rect 1562 22953 1597 22987
rect 1631 22953 1666 22987
rect 1700 22953 1735 22987
rect 1769 22953 1804 22987
rect 1838 22953 1873 22987
rect 1907 22953 1942 22987
rect 1976 22953 2011 22987
rect 2045 22953 2080 22987
rect 2114 22953 2149 22987
rect 1286 22919 2149 22953
rect 1286 22885 1321 22919
rect 1355 22885 1390 22919
rect 1424 22885 1459 22919
rect 1493 22885 1528 22919
rect 1562 22885 1597 22919
rect 1631 22885 1666 22919
rect 1700 22885 1735 22919
rect 1769 22885 1804 22919
rect 1838 22885 1873 22919
rect 1907 22885 1942 22919
rect 1976 22885 2011 22919
rect 2045 22885 2080 22919
rect 2114 22885 2149 22919
rect 776 22850 912 22885
rect 810 22816 844 22850
rect 878 22817 912 22850
rect 1286 22851 2149 22885
rect 1286 22817 1321 22851
rect 1355 22817 1390 22851
rect 1424 22817 1459 22851
rect 1493 22817 1528 22851
rect 1562 22817 1597 22851
rect 1631 22817 1666 22851
rect 1700 22817 1735 22851
rect 1769 22817 1804 22851
rect 1838 22817 1873 22851
rect 1907 22817 1942 22851
rect 1976 22817 2011 22851
rect 2045 22817 2080 22851
rect 2114 22817 2149 22851
rect 878 22816 946 22817
rect 776 22782 946 22816
rect 776 22781 912 22782
rect 810 22747 844 22781
rect 878 22748 912 22781
rect 878 22747 946 22748
rect 776 22713 946 22747
rect 776 22712 912 22713
rect 810 22678 844 22712
rect 878 22679 912 22712
rect 878 22678 946 22679
rect 776 22644 946 22678
rect 776 22643 912 22644
rect 810 22609 844 22643
rect 878 22610 912 22643
rect 878 22609 946 22610
rect 776 22575 946 22609
rect 776 22574 912 22575
rect 810 22540 844 22574
rect 878 22541 912 22574
rect 878 22540 946 22541
rect 776 22506 946 22540
rect 776 22505 912 22506
rect 810 22471 844 22505
rect 878 22472 912 22505
rect 878 22471 946 22472
rect 776 22437 946 22471
rect 776 22436 912 22437
rect 810 22402 844 22436
rect 878 22403 912 22436
rect 878 22402 946 22403
rect 776 22368 946 22402
rect 776 22367 912 22368
rect 810 22333 844 22367
rect 878 22334 912 22367
rect 878 22333 946 22334
rect 776 22299 946 22333
rect 776 22298 912 22299
rect 810 22264 844 22298
rect 878 22265 912 22298
rect 878 22264 946 22265
rect 776 22230 946 22264
rect 776 22229 912 22230
rect 810 22195 844 22229
rect 878 22196 912 22229
rect 878 22195 946 22196
rect 776 22161 946 22195
rect 776 22160 912 22161
rect 810 22126 844 22160
rect 878 22127 912 22160
rect 878 22126 946 22127
rect 776 22092 946 22126
rect 776 22091 912 22092
rect 810 22057 844 22091
rect 878 22058 912 22091
rect 878 22057 946 22058
rect 776 22023 946 22057
rect 776 22022 912 22023
rect 810 21988 844 22022
rect 878 21989 912 22022
rect 878 21988 946 21989
rect 776 21954 946 21988
rect 776 21953 912 21954
rect 810 21919 844 21953
rect 878 21920 912 21953
rect 878 21919 946 21920
rect 776 21885 946 21919
rect 776 21884 912 21885
rect 810 21850 844 21884
rect 878 21851 912 21884
rect 878 21850 946 21851
rect 776 21816 946 21850
rect 776 21815 912 21816
rect 810 21781 844 21815
rect 878 21782 912 21815
rect 878 21781 946 21782
rect 776 21747 946 21781
rect 776 21746 912 21747
rect 810 21712 844 21746
rect 878 21713 912 21746
rect 878 21712 946 21713
rect 776 21678 946 21712
rect 776 21677 912 21678
rect 810 21643 844 21677
rect 878 21644 912 21677
rect 878 21643 946 21644
rect 776 21609 946 21643
rect 776 21608 912 21609
rect 810 21574 844 21608
rect 878 21575 912 21608
rect 878 21574 946 21575
rect 776 21540 946 21574
rect 776 21539 912 21540
rect 810 21505 844 21539
rect 878 21506 912 21539
rect 878 21505 946 21506
rect 776 21471 946 21505
rect 776 21470 912 21471
rect 810 21436 844 21470
rect 878 21437 912 21470
rect 878 21436 946 21437
rect 776 21402 946 21436
rect 776 21401 912 21402
rect 810 21367 844 21401
rect 878 21368 912 21401
rect 878 21367 946 21368
rect 776 21333 946 21367
rect 776 21332 912 21333
rect 810 21298 844 21332
rect 878 21299 912 21332
rect 878 21298 946 21299
rect 776 21264 946 21298
rect 776 21263 912 21264
rect 810 21229 844 21263
rect 878 21230 912 21263
rect 878 21229 946 21230
rect 776 21195 946 21229
rect 776 21194 912 21195
rect 810 21160 844 21194
rect 878 21161 912 21194
rect 878 21160 946 21161
rect 776 21126 946 21160
rect 776 21125 912 21126
rect 810 21091 844 21125
rect 878 21092 912 21125
rect 878 21091 946 21092
rect 776 21057 946 21091
rect 776 21056 912 21057
rect 810 21022 844 21056
rect 878 21023 912 21056
rect 878 21022 946 21023
rect 776 20988 946 21022
rect 776 20987 912 20988
rect 810 20953 844 20987
rect 878 20954 912 20987
rect 878 20953 946 20954
rect 776 20919 946 20953
rect 776 20918 912 20919
rect 810 20884 844 20918
rect 878 20885 912 20918
rect 878 20884 946 20885
rect 776 20850 946 20884
rect 776 20849 912 20850
rect 810 20815 844 20849
rect 878 20816 912 20849
rect 878 20815 946 20816
rect 776 20781 946 20815
rect 776 20780 912 20781
rect 810 20746 844 20780
rect 878 20747 912 20780
rect 878 20746 946 20747
rect 776 20712 946 20746
rect 776 20711 912 20712
rect 810 20677 844 20711
rect 878 20678 912 20711
rect 878 20677 946 20678
rect 776 20643 946 20677
rect 776 20642 912 20643
rect 810 20608 844 20642
rect 878 20609 912 20642
rect 878 20608 946 20609
rect 776 20574 946 20608
rect 776 20573 912 20574
rect 810 20539 844 20573
rect 878 20540 912 20573
rect 878 20539 946 20540
rect 776 20505 946 20539
rect 776 20504 912 20505
rect 810 20470 844 20504
rect 878 20471 912 20504
rect 878 20470 946 20471
rect 776 20436 946 20470
rect 776 20435 912 20436
rect 810 20401 844 20435
rect 878 20402 912 20435
rect 878 20401 946 20402
rect 776 20367 946 20401
rect 776 20366 912 20367
rect 810 20332 844 20366
rect 878 20333 912 20366
rect 878 20332 946 20333
rect 776 20298 946 20332
rect 776 20297 912 20298
rect 810 20263 844 20297
rect 878 20264 912 20297
rect 878 20263 946 20264
rect 776 20229 946 20263
rect 776 20228 912 20229
rect 810 20194 844 20228
rect 878 20195 912 20228
rect 878 20194 946 20195
rect 776 20160 946 20194
rect 776 20159 912 20160
rect 810 20125 844 20159
rect 878 20126 912 20159
rect 878 20125 946 20126
rect 776 20091 946 20125
rect 776 20090 912 20091
rect 810 20056 844 20090
rect 878 20057 912 20090
rect 878 20056 946 20057
rect 776 20022 946 20056
rect 776 20021 912 20022
rect 810 19987 844 20021
rect 878 19988 912 20021
rect 878 19987 946 19988
rect 776 19953 946 19987
rect 776 19952 912 19953
rect 810 19918 844 19952
rect 878 19919 912 19952
rect 878 19918 946 19919
rect 776 19884 946 19918
rect 776 19883 912 19884
rect 810 19849 844 19883
rect 878 19850 912 19883
rect 878 19849 946 19850
rect 776 19815 946 19849
rect 776 19814 912 19815
rect 810 19780 844 19814
rect 878 19781 912 19814
rect 878 19780 946 19781
rect 776 19746 946 19780
rect 776 19745 912 19746
rect 810 19711 844 19745
rect 878 19712 912 19745
rect 878 19711 946 19712
rect 776 19677 946 19711
rect 776 19676 912 19677
rect 810 19642 844 19676
rect 878 19643 912 19676
rect 878 19642 946 19643
rect 776 19608 946 19642
rect 776 19607 912 19608
rect 810 19573 844 19607
rect 878 19574 912 19607
rect 878 19573 946 19574
rect 776 19539 946 19573
rect 776 19538 912 19539
rect 810 19504 844 19538
rect 878 19505 912 19538
rect 878 19504 946 19505
rect 776 19470 946 19504
rect 776 19469 912 19470
rect 810 19435 844 19469
rect 878 19436 912 19469
rect 878 19435 946 19436
rect 776 19401 946 19435
rect 776 19400 912 19401
rect 810 19366 844 19400
rect 878 19367 912 19400
rect 878 19366 946 19367
rect 776 19332 946 19366
rect 776 19331 912 19332
rect 810 19297 844 19331
rect 878 19298 912 19331
rect 878 19297 946 19298
rect 776 19263 946 19297
rect 776 19262 912 19263
rect 810 19228 844 19262
rect 878 19229 912 19262
rect 878 19228 946 19229
rect 776 19194 946 19228
rect 776 19193 912 19194
rect 810 19159 844 19193
rect 878 19160 912 19193
rect 878 19159 946 19160
rect 776 19125 946 19159
rect 776 19124 912 19125
rect 810 19090 844 19124
rect 878 19091 912 19124
rect 878 19090 946 19091
rect 776 19056 946 19090
rect 776 19055 912 19056
rect 810 19021 844 19055
rect 878 19022 912 19055
rect 878 19021 946 19022
rect 776 18987 946 19021
rect 776 18986 912 18987
rect 810 18952 844 18986
rect 878 18953 912 18986
rect 878 18952 946 18953
rect 776 18918 946 18952
rect 776 18917 912 18918
rect 810 18883 844 18917
rect 878 18884 912 18917
rect 878 18883 946 18884
rect 776 18849 946 18883
rect 776 18848 912 18849
rect 810 18814 844 18848
rect 878 18815 912 18848
rect 878 18814 946 18815
rect 776 18780 946 18814
rect 776 18779 912 18780
rect 810 18745 844 18779
rect 878 18746 912 18779
rect 878 18745 946 18746
rect 776 18711 946 18745
rect 776 18710 912 18711
rect 810 18676 844 18710
rect 878 18677 912 18710
rect 878 18676 946 18677
rect 776 18642 946 18676
rect 776 18641 912 18642
rect 810 18607 844 18641
rect 878 18608 912 18641
rect 878 18607 946 18608
rect 776 18573 946 18607
rect 776 18572 912 18573
rect 810 18538 844 18572
rect 878 18539 912 18572
rect 878 18538 946 18539
rect 776 18504 946 18538
rect 776 18503 912 18504
rect 810 18469 844 18503
rect 878 18470 912 18503
rect 878 18469 946 18470
rect 776 18435 946 18469
rect 776 18434 912 18435
rect 810 18400 844 18434
rect 878 18401 912 18434
rect 878 18400 946 18401
rect 776 18366 946 18400
rect 776 18365 912 18366
rect 878 18332 912 18365
rect 878 18297 946 18332
rect 1090 22667 1832 22673
rect 1090 22631 1174 22667
rect 1208 22633 1252 22667
rect 1286 22665 1330 22667
rect 1364 22665 1408 22667
rect 1442 22665 1486 22667
rect 1520 22665 1564 22667
rect 1598 22665 1642 22667
rect 1676 22665 1720 22667
rect 1754 22665 1832 22667
rect 1286 22633 1314 22665
rect 1208 22631 1314 22633
rect 1090 22597 1314 22631
rect 1090 22595 1098 22597
rect 1200 22595 1314 22597
rect 1756 22595 1832 22665
rect 1090 22561 1096 22595
rect 1202 22561 1252 22595
rect 1286 22563 1314 22595
rect 1286 22561 1330 22563
rect 1364 22561 1408 22563
rect 1442 22561 1486 22563
rect 1520 22561 1564 22563
rect 1598 22561 1642 22563
rect 1676 22561 1720 22563
rect 1090 22522 1098 22561
rect 1200 22555 1720 22561
rect 1200 22522 1208 22555
rect 1090 22488 1096 22522
rect 1202 22488 1208 22522
rect 1090 22449 1098 22488
rect 1200 22449 1208 22488
rect 1090 22415 1096 22449
rect 1202 22415 1208 22449
rect 1090 22376 1098 22415
rect 1200 22376 1208 22415
rect 1714 22489 1720 22555
rect 1826 22489 1832 22595
rect 1714 22450 1722 22489
rect 1824 22450 1832 22489
rect 1714 22416 1720 22450
rect 1826 22416 1832 22450
rect 1090 22342 1096 22376
rect 1202 22342 1208 22376
rect 1350 22404 1417 22411
rect 1350 22363 1366 22404
rect 1090 22303 1098 22342
rect 1200 22303 1208 22342
rect 1090 22269 1096 22303
rect 1202 22269 1208 22303
rect 1400 22363 1417 22404
rect 1506 22404 1573 22411
rect 1506 22363 1522 22404
rect 1366 22321 1400 22359
rect 1556 22363 1573 22404
rect 1714 22377 1722 22416
rect 1824 22377 1832 22416
rect 1522 22321 1556 22359
rect 1714 22343 1720 22377
rect 1826 22343 1832 22377
rect 1714 22304 1722 22343
rect 1824 22304 1832 22343
rect 1090 22230 1098 22269
rect 1200 22230 1208 22269
rect 1714 22270 1720 22304
rect 1826 22270 1832 22304
rect 1090 22196 1096 22230
rect 1202 22196 1208 22230
rect 1090 22157 1098 22196
rect 1200 22157 1208 22196
rect 1090 22123 1096 22157
rect 1202 22123 1208 22157
rect 1090 22084 1098 22123
rect 1200 22084 1208 22123
rect 1090 22050 1096 22084
rect 1202 22050 1208 22084
rect 1090 22011 1098 22050
rect 1200 22011 1208 22050
rect 1090 21977 1096 22011
rect 1202 21977 1208 22011
rect 1090 21938 1098 21977
rect 1200 21938 1208 21977
rect 1090 16432 1096 21938
rect 1202 16472 1208 21938
rect 1288 22255 1322 22259
rect 1288 22183 1322 22209
rect 1288 22111 1322 22141
rect 1288 22039 1322 22073
rect 1288 21971 1322 22005
rect 1288 21903 1322 21933
rect 1288 21835 1322 21861
rect 1288 21767 1322 21789
rect 1444 22255 1478 22259
rect 1444 22183 1478 22209
rect 1444 22111 1478 22141
rect 1444 22039 1478 22073
rect 1444 21971 1478 22005
rect 1444 21903 1478 21933
rect 1444 21835 1478 21861
rect 1444 21767 1478 21789
rect 1600 22255 1634 22259
rect 1600 22183 1634 22209
rect 1600 22111 1634 22141
rect 1600 22039 1634 22073
rect 1600 21971 1634 22005
rect 1600 21903 1634 21933
rect 1600 21835 1634 21861
rect 1600 21767 1634 21789
rect 1714 22231 1722 22270
rect 1824 22231 1832 22270
rect 1714 22197 1720 22231
rect 1826 22197 1832 22231
rect 1714 22158 1722 22197
rect 1824 22158 1832 22197
rect 1714 22124 1720 22158
rect 1826 22124 1832 22158
rect 1714 22085 1722 22124
rect 1824 22085 1832 22124
rect 1714 22051 1720 22085
rect 1826 22051 1832 22085
rect 1714 22012 1722 22051
rect 1824 22012 1832 22051
rect 1714 21978 1720 22012
rect 1826 21978 1832 22012
rect 1714 21939 1722 21978
rect 1824 21939 1832 21978
rect 1714 21905 1720 21939
rect 1826 21905 1832 21939
rect 1714 21866 1722 21905
rect 1824 21866 1832 21905
rect 1714 21832 1720 21866
rect 1826 21832 1832 21866
rect 1714 21793 1722 21832
rect 1824 21793 1832 21832
rect 1714 21759 1720 21793
rect 1826 21759 1832 21793
rect 1714 21720 1722 21759
rect 1824 21720 1832 21759
rect 1350 21674 1366 21679
rect 1400 21674 1417 21679
rect 1350 21672 1417 21674
rect 1350 21638 1366 21672
rect 1400 21638 1417 21672
rect 1350 21636 1417 21638
rect 1350 21631 1366 21636
rect 1400 21631 1417 21636
rect 1506 21674 1522 21679
rect 1714 21686 1720 21720
rect 1826 21686 1832 21720
rect 1556 21674 1573 21679
rect 1506 21672 1573 21674
rect 1506 21638 1522 21672
rect 1556 21638 1573 21672
rect 1506 21636 1573 21638
rect 1506 21631 1522 21636
rect 1556 21631 1573 21636
rect 1714 21647 1722 21686
rect 1824 21647 1832 21686
rect 1714 21613 1720 21647
rect 1826 21613 1832 21647
rect 1288 21521 1322 21543
rect 1288 21449 1322 21475
rect 1288 21377 1322 21407
rect 1288 21305 1322 21339
rect 1288 21237 1322 21271
rect 1288 21169 1322 21199
rect 1288 21101 1322 21127
rect 1288 21051 1322 21055
rect 1444 21521 1478 21543
rect 1444 21449 1478 21475
rect 1444 21377 1478 21407
rect 1444 21305 1478 21339
rect 1444 21237 1478 21271
rect 1444 21169 1478 21199
rect 1444 21101 1478 21127
rect 1444 21051 1478 21055
rect 1600 21521 1634 21543
rect 1600 21449 1634 21475
rect 1600 21377 1634 21407
rect 1600 21305 1634 21339
rect 1600 21237 1634 21271
rect 1600 21169 1634 21199
rect 1600 21101 1634 21127
rect 1714 21574 1722 21613
rect 1824 21574 1832 21613
rect 1714 21540 1720 21574
rect 1826 21540 1832 21574
rect 1714 21501 1722 21540
rect 1824 21501 1832 21540
rect 1714 21467 1720 21501
rect 1826 21467 1832 21501
rect 1714 21428 1722 21467
rect 1824 21428 1832 21467
rect 1714 21394 1720 21428
rect 1826 21394 1832 21428
rect 1714 21355 1722 21394
rect 1824 21355 1832 21394
rect 1714 21321 1720 21355
rect 1826 21321 1832 21355
rect 1714 21282 1722 21321
rect 1824 21282 1832 21321
rect 1714 21248 1720 21282
rect 1826 21248 1832 21282
rect 1714 21209 1722 21248
rect 1824 21209 1832 21248
rect 1714 21175 1720 21209
rect 1826 21175 1832 21209
rect 1714 21136 1722 21175
rect 1824 21136 1832 21175
rect 1714 21102 1720 21136
rect 1826 21102 1832 21136
rect 1714 21070 1722 21102
rect 1600 21051 1634 21055
rect 1824 21070 1832 21102
rect 1714 16472 1722 16473
rect 1202 16466 1722 16472
rect 1202 16464 1244 16466
rect 1278 16464 1320 16466
rect 1354 16464 1395 16466
rect 1429 16464 1470 16466
rect 1504 16464 1545 16466
rect 1579 16464 1620 16466
rect 1654 16464 1695 16466
rect 1676 16432 1695 16464
rect 1090 16362 1166 16432
rect 1676 16430 1722 16432
rect 1824 16430 1832 16473
rect 1676 16417 1832 16430
rect 1676 16396 1792 16417
rect 1676 16362 1710 16396
rect 1744 16394 1792 16396
rect 1748 16383 1792 16394
rect 1826 16383 1832 16417
rect 1090 16360 1168 16362
rect 1202 16360 1246 16362
rect 1280 16360 1324 16362
rect 1358 16360 1402 16362
rect 1436 16360 1480 16362
rect 1514 16360 1558 16362
rect 1592 16360 1636 16362
rect 1670 16360 1714 16362
rect 1748 16360 1832 16383
rect 1090 16354 1832 16360
rect 2217 16418 2387 16453
rect 2251 16384 2285 16418
rect 2319 16384 2353 16418
rect 2217 16349 2387 16384
rect 2251 16315 2285 16349
rect 2319 16315 2353 16349
rect 2217 16280 2387 16315
rect 2251 16246 2285 16280
rect 2319 16246 2353 16280
rect 2217 16211 2387 16246
rect 946 16155 981 16189
rect 1015 16155 1050 16189
rect 1084 16155 1119 16189
rect 1153 16155 1188 16189
rect 1222 16155 1257 16189
rect 1291 16155 1326 16189
rect 1360 16155 1395 16189
rect 1429 16155 1464 16189
rect 1498 16155 1533 16189
rect 1567 16155 1602 16189
rect 1636 16155 1671 16189
rect 1705 16155 1740 16189
rect 1774 16155 1809 16189
rect 878 16121 1809 16155
rect 2183 16177 2217 16189
rect 2251 16177 2285 16211
rect 2319 16177 2353 16211
rect 2183 16142 2387 16177
rect 878 16087 913 16121
rect 947 16087 982 16121
rect 1016 16087 1051 16121
rect 1085 16087 1120 16121
rect 1154 16087 1189 16121
rect 1223 16087 1258 16121
rect 1292 16087 1327 16121
rect 1361 16087 1396 16121
rect 1430 16087 1465 16121
rect 1499 16087 1534 16121
rect 1568 16087 1603 16121
rect 1637 16087 1672 16121
rect 1706 16087 1741 16121
rect 776 16053 1741 16087
rect 776 16019 844 16053
rect 878 16019 913 16053
rect 947 16019 982 16053
rect 1016 16019 1051 16053
rect 1085 16019 1120 16053
rect 1154 16019 1189 16053
rect 1223 16019 1258 16053
rect 1292 16019 1327 16053
rect 1361 16019 1396 16053
rect 1430 16019 1465 16053
rect 1499 16019 1534 16053
rect 1568 16019 1603 16053
rect 1637 16019 1672 16053
rect 1706 16019 1741 16053
rect 2183 16108 2217 16142
rect 2251 16108 2285 16142
rect 2319 16108 2353 16142
rect 2183 16073 2387 16108
rect 2183 16039 2217 16073
rect 2251 16039 2285 16073
rect 2319 16039 2353 16073
rect 2183 16019 2387 16039
rect 2217 16004 2387 16019
rect 2251 15970 2285 16004
rect 2319 15970 2353 16004
rect 2217 15935 2387 15970
rect 2251 15901 2285 15935
rect 2319 15901 2353 15935
rect 2217 15866 2387 15901
rect 2251 15832 2285 15866
rect 2319 15832 2353 15866
rect 2217 15797 2387 15832
rect 2251 15763 2285 15797
rect 2319 15763 2353 15797
rect 2217 15728 2387 15763
rect 2251 15694 2285 15728
rect 2319 15694 2353 15728
rect 2217 15659 2387 15694
rect 2251 15625 2285 15659
rect 2319 15625 2353 15659
rect 2217 15591 2387 15625
rect 69 13625 192 13659
rect 226 13625 260 13659
rect 69 13591 260 13625
rect 171 13557 260 13591
rect 171 13523 328 13557
rect 239 13489 328 13523
rect 26678 13489 26712 13659
rect 26627 13415 26797 13489
rect 507 13226 26404 13232
rect 507 13154 585 13226
rect 619 13222 658 13226
rect 692 13222 731 13226
rect 765 13222 804 13226
rect 507 9736 513 13154
rect 26326 13154 26404 13226
rect 26398 13120 26404 13154
rect 619 13082 653 13120
rect 26254 13086 26292 13120
rect 691 13048 730 13052
rect 764 13048 803 13052
rect 837 13048 876 13052
rect 26394 13080 26404 13120
rect 691 13042 26224 13048
rect 26398 13046 26404 13080
rect 691 9808 697 13042
rect 26214 13008 26224 13042
rect 26214 12974 26220 13008
rect 26394 13006 26404 13046
rect 26214 12934 26224 12974
rect 26398 12972 26404 13006
rect 26214 12900 26220 12934
rect 26394 12932 26404 12972
rect 26214 12860 26224 12900
rect 26398 12898 26404 12932
rect 619 9769 697 9808
rect 619 9748 657 9769
rect 507 9714 517 9736
rect 551 9714 585 9736
rect 619 9714 653 9748
rect 691 9735 697 9769
rect 687 9714 697 9735
rect 507 9697 697 9714
rect 507 9663 513 9697
rect 547 9679 585 9697
rect 619 9696 697 9697
rect 619 9679 657 9696
rect 507 9645 517 9663
rect 551 9645 585 9679
rect 619 9645 653 9679
rect 691 9662 697 9696
rect 687 9645 697 9662
rect 507 9624 697 9645
rect 507 9590 513 9624
rect 547 9610 585 9624
rect 619 9623 697 9624
rect 619 9610 657 9623
rect 507 9576 517 9590
rect 551 9576 585 9610
rect 619 9576 653 9610
rect 691 9589 697 9623
rect 687 9576 697 9589
rect 507 9551 697 9576
rect 507 9517 513 9551
rect 547 9541 585 9551
rect 619 9550 697 9551
rect 619 9541 657 9550
rect 507 9507 517 9517
rect 551 9507 585 9541
rect 619 9507 653 9541
rect 691 9516 697 9550
rect 687 9507 697 9516
rect 507 9478 697 9507
rect 507 9444 513 9478
rect 547 9472 585 9478
rect 619 9477 697 9478
rect 619 9472 657 9477
rect 507 9438 517 9444
rect 551 9438 585 9472
rect 619 9438 653 9472
rect 691 9443 697 9477
rect 687 9438 697 9443
rect 507 9405 697 9438
rect 507 9371 513 9405
rect 547 9403 585 9405
rect 619 9404 697 9405
rect 619 9403 657 9404
rect 507 9369 517 9371
rect 551 9369 585 9403
rect 619 9369 653 9403
rect 691 9370 697 9404
rect 687 9369 697 9370
rect 507 9334 697 9369
rect 507 9332 517 9334
rect 507 9298 513 9332
rect 551 9300 585 9334
rect 619 9300 653 9334
rect 687 9331 697 9334
rect 547 9298 585 9300
rect 619 9298 657 9300
rect 507 9297 657 9298
rect 691 9297 697 9331
rect 507 9265 697 9297
rect 507 9259 517 9265
rect 507 9225 513 9259
rect 551 9231 585 9265
rect 619 9231 653 9265
rect 687 9258 697 9265
rect 547 9225 585 9231
rect 619 9225 657 9231
rect 507 9224 657 9225
rect 691 9224 697 9258
rect 507 9196 697 9224
rect 507 9186 517 9196
rect 507 9152 513 9186
rect 551 9162 585 9196
rect 619 9162 653 9196
rect 687 9185 697 9196
rect 547 9152 585 9162
rect 619 9152 657 9162
rect 507 9151 657 9152
rect 691 9151 697 9185
rect 507 9127 697 9151
rect 507 9113 517 9127
rect 507 9079 513 9113
rect 551 9093 585 9127
rect 619 9093 653 9127
rect 687 9112 697 9127
rect 547 9079 585 9093
rect 619 9079 657 9093
rect 507 9078 657 9079
rect 691 9078 697 9112
rect 507 9058 697 9078
rect 507 9040 517 9058
rect 507 9006 513 9040
rect 551 9024 585 9058
rect 619 9024 653 9058
rect 687 9039 697 9058
rect 547 9006 585 9024
rect 619 9006 657 9024
rect 507 9005 657 9006
rect 691 9005 697 9039
rect 507 8989 697 9005
rect 507 8967 517 8989
rect 507 8933 513 8967
rect 551 8955 585 8989
rect 619 8955 653 8989
rect 687 8966 697 8989
rect 547 8933 585 8955
rect 619 8933 657 8955
rect 507 8932 657 8933
rect 691 8932 697 8966
rect 507 8920 697 8932
rect 507 8894 517 8920
rect 507 8860 513 8894
rect 551 8886 585 8920
rect 619 8886 653 8920
rect 687 8893 697 8920
rect 547 8860 585 8886
rect 619 8860 657 8886
rect 507 8859 657 8860
rect 691 8859 697 8893
rect 507 8851 697 8859
rect 507 8821 517 8851
rect 507 8787 513 8821
rect 551 8817 585 8851
rect 619 8817 653 8851
rect 687 8820 697 8851
rect 547 8787 585 8817
rect 619 8787 657 8817
rect 507 8786 657 8787
rect 691 8786 697 8820
rect 507 8782 697 8786
rect 507 8748 517 8782
rect 551 8748 585 8782
rect 619 8748 653 8782
rect 687 8748 697 8782
rect 507 8714 513 8748
rect 547 8714 585 8748
rect 619 8747 697 8748
rect 619 8714 657 8747
rect 507 8713 657 8714
rect 691 8713 697 8747
rect 507 8679 517 8713
rect 551 8679 585 8713
rect 619 8679 653 8713
rect 687 8679 697 8713
rect 507 8675 697 8679
rect 507 8641 513 8675
rect 547 8644 585 8675
rect 619 8674 697 8675
rect 619 8644 657 8674
rect 507 8610 517 8641
rect 551 8610 585 8644
rect 619 8610 653 8644
rect 691 8640 697 8674
rect 687 8610 697 8640
rect 507 8602 697 8610
rect 507 8568 513 8602
rect 547 8575 585 8602
rect 619 8601 697 8602
rect 619 8575 657 8601
rect 507 8541 517 8568
rect 551 8541 585 8575
rect 619 8541 653 8575
rect 691 8567 697 8601
rect 687 8541 697 8567
rect 507 8529 697 8541
rect 507 8495 513 8529
rect 547 8506 585 8529
rect 619 8528 697 8529
rect 619 8506 657 8528
rect 507 8472 517 8495
rect 551 8472 585 8506
rect 619 8472 653 8506
rect 691 8494 697 8528
rect 687 8472 697 8494
rect 507 8456 697 8472
rect 507 8422 513 8456
rect 547 8437 585 8456
rect 619 8455 697 8456
rect 619 8437 657 8455
rect 507 8403 517 8422
rect 551 8403 585 8437
rect 619 8403 653 8437
rect 691 8421 697 8455
rect 687 8403 697 8421
rect 507 8383 697 8403
rect 507 8349 513 8383
rect 547 8368 585 8383
rect 619 8382 697 8383
rect 619 8368 657 8382
rect 507 8334 517 8349
rect 551 8334 585 8368
rect 619 8334 653 8368
rect 691 8348 697 8382
rect 687 8334 697 8348
rect 507 8310 697 8334
rect 507 8276 513 8310
rect 547 8299 585 8310
rect 619 8309 697 8310
rect 619 8299 657 8309
rect 507 8237 517 8276
rect 691 8275 697 8309
rect 507 8203 513 8237
rect 687 8236 697 8275
rect 507 8164 517 8203
rect 691 8202 697 8236
rect 507 8130 513 8164
rect 687 8163 697 8202
rect 507 8091 517 8130
rect 691 8129 697 8163
rect 507 8057 513 8091
rect 687 8090 697 8129
rect 507 8018 517 8057
rect 691 8056 697 8090
rect 507 7984 513 8018
rect 687 8017 697 8056
rect 507 7945 517 7984
rect 691 7983 697 8017
rect 507 7911 513 7945
rect 687 7944 697 7983
rect 507 7872 517 7911
rect 691 7910 697 7944
rect 507 7838 513 7872
rect 687 7871 697 7910
rect 507 7799 517 7838
rect 691 7837 697 7871
rect 507 7765 513 7799
rect 687 7798 697 7837
rect 507 7726 517 7765
rect 691 7764 697 7798
rect 507 7692 513 7726
rect 687 7725 697 7764
rect 507 7653 517 7692
rect 691 7691 697 7725
rect 507 7619 513 7653
rect 687 7652 697 7691
rect 507 7580 517 7619
rect 691 7618 697 7652
rect 507 7546 513 7580
rect 687 7579 697 7618
rect 507 7507 517 7546
rect 691 7545 697 7579
rect 507 7473 513 7507
rect 687 7506 697 7545
rect 507 7434 517 7473
rect 691 7472 697 7506
rect 507 7400 513 7434
rect 687 7433 697 7472
rect 507 7361 517 7400
rect 691 7399 697 7433
rect 507 7327 513 7361
rect 687 7360 697 7399
rect 507 7288 517 7327
rect 691 7326 697 7360
rect 507 7254 513 7288
rect 687 7287 697 7326
rect 507 7215 517 7254
rect 691 7253 697 7287
rect 507 7181 513 7215
rect 687 7214 697 7253
rect 507 7142 517 7181
rect 691 7180 697 7214
rect 507 7108 513 7142
rect 687 7141 697 7180
rect 507 7069 517 7108
rect 691 7107 697 7141
rect 507 7035 513 7069
rect 687 7068 697 7107
rect 507 6996 517 7035
rect 691 7034 697 7068
rect 507 6962 513 6996
rect 687 6995 697 7034
rect 507 6923 517 6962
rect 691 6961 697 6995
rect 507 6889 513 6923
rect 687 6922 697 6961
rect 507 6850 517 6889
rect 691 6888 697 6922
rect 507 6816 513 6850
rect 687 6849 697 6888
rect 507 6777 517 6816
rect 691 6815 697 6849
rect 507 6743 513 6777
rect 687 6776 697 6815
rect 507 6704 517 6743
rect 691 6742 697 6776
rect 507 6670 513 6704
rect 687 6703 697 6742
rect 507 6631 517 6670
rect 691 6669 697 6703
rect 507 6597 513 6631
rect 687 6630 697 6669
rect 893 12840 26006 12846
rect 893 12806 971 12840
rect 1005 12837 1044 12840
rect 1078 12837 1117 12840
rect 1151 12837 1190 12840
rect 1224 12837 1263 12840
rect 1297 12837 1336 12840
rect 1370 12837 1409 12840
rect 1443 12837 1482 12840
rect 1516 12837 1555 12840
rect 1589 12837 1628 12840
rect 1662 12837 1701 12840
rect 1735 12837 1774 12840
rect 1019 12806 1044 12837
rect 893 12803 985 12806
rect 1019 12803 1053 12806
rect 893 12769 1053 12803
rect 893 12768 903 12769
rect 1005 12768 1053 12769
rect 893 9638 899 12768
rect 1005 12734 1044 12768
rect 1078 12734 1117 12735
rect 25928 12768 26006 12840
rect 25928 12736 25966 12768
rect 25928 12734 25941 12736
rect 26000 12734 26006 12768
rect 1005 12701 1121 12734
rect 1073 12696 1121 12701
rect 1077 12662 1116 12696
rect 25856 12702 25941 12734
rect 25975 12702 26006 12734
rect 25856 12694 26006 12702
rect 25856 12668 25894 12694
rect 25928 12668 25966 12694
rect 1150 12662 1189 12667
rect 1223 12662 1262 12667
rect 1296 12662 1335 12667
rect 1369 12662 1408 12667
rect 1442 12662 1481 12667
rect 1515 12662 1554 12667
rect 1588 12662 1627 12667
rect 1661 12662 1700 12667
rect 1734 12662 1773 12667
rect 1807 12662 1846 12667
rect 25856 12662 25873 12668
rect 1077 12656 25873 12662
rect 26000 12660 26006 12694
rect 1077 9710 1083 12656
rect 25805 12622 25873 12656
rect 25805 12600 25822 12622
rect 25856 12600 25873 12622
rect 25975 12620 26006 12660
rect 26000 12586 26006 12620
rect 25975 12546 26006 12586
rect 26000 12512 26006 12546
rect 25975 12472 26006 12512
rect 26000 12438 26006 12472
rect 25975 12398 26006 12438
rect 26000 12364 26006 12398
rect 25975 12325 26006 12364
rect 26000 12291 26006 12325
rect 25975 12252 26006 12291
rect 26000 12218 26006 12252
rect 25975 12142 26006 12218
rect 26000 12108 26006 12142
rect 25975 12069 26006 12108
rect 26000 12035 26006 12069
rect 25975 11996 26006 12035
rect 26000 11962 26006 11996
rect 25975 11923 26006 11962
rect 26000 11889 26006 11923
rect 25975 11850 26006 11889
rect 26000 11816 26006 11850
rect 25975 11777 26006 11816
rect 26000 11743 26006 11777
rect 25975 11704 26006 11743
rect 26000 11670 26006 11704
rect 25975 11631 26006 11670
rect 26000 11597 26006 11631
rect 25975 11558 26006 11597
rect 26000 11524 26006 11558
rect 25975 11485 26006 11524
rect 26000 11451 26006 11485
rect 25975 11412 26006 11451
rect 26000 11378 26006 11412
rect 25975 11339 26006 11378
rect 26000 11305 26006 11339
rect 25975 11266 26006 11305
rect 26000 11232 26006 11266
rect 25975 11193 26006 11232
rect 26000 11159 26006 11193
rect 25975 11120 26006 11159
rect 26000 11086 26006 11120
rect 25975 11047 26006 11086
rect 26000 11013 26006 11047
rect 25975 10974 26006 11013
rect 26000 10940 26006 10974
rect 25975 10901 26006 10940
rect 26000 10867 26006 10901
rect 25975 10828 26006 10867
rect 26000 10794 26006 10828
rect 25975 10755 26006 10794
rect 26000 10721 26006 10755
rect 25975 10682 26006 10721
rect 26000 10648 26006 10682
rect 25975 10609 26006 10648
rect 1732 10584 1988 10591
rect 1335 10550 1382 10584
rect 1416 10550 1462 10584
rect 1496 10550 1542 10584
rect 1576 10550 1622 10584
rect 1656 10550 1702 10584
rect 1736 10550 1748 10584
rect 1816 10550 1843 10584
rect 1896 10550 1938 10584
rect 1976 10550 1988 10584
rect 1732 10543 1988 10550
rect 26000 10575 26006 10609
rect 25975 10536 26006 10575
rect 26000 10502 26006 10536
rect 1687 10426 1721 10449
rect 1687 10352 1721 10381
rect 1687 10279 1721 10313
rect 1687 10211 1721 10245
rect 1687 10143 1721 10177
rect 1687 10075 1721 10109
rect 1687 10007 1721 10041
rect 1687 9957 1721 9973
rect 1843 10483 1877 10499
rect 1843 10415 1877 10449
rect 1843 10347 1877 10381
rect 1843 10279 1877 10313
rect 1843 10211 1877 10245
rect 1843 10149 1877 10177
rect 1843 10077 1877 10109
rect 1843 10007 1877 10041
rect 1843 9957 1877 9973
rect 1999 10426 2033 10449
rect 1999 10352 2033 10381
rect 1999 10279 2033 10313
rect 1999 10211 2033 10245
rect 1999 10143 2033 10177
rect 1999 10075 2033 10109
rect 1999 10007 2033 10041
rect 1999 9957 2033 9973
rect 25975 10463 26006 10502
rect 26000 10429 26006 10463
rect 25975 10390 26006 10429
rect 26000 10356 26006 10390
rect 25975 10317 26006 10356
rect 26000 10283 26006 10317
rect 25975 10244 26006 10283
rect 26000 10210 26006 10244
rect 25975 10171 26006 10210
rect 26000 10137 26006 10171
rect 25975 10098 26006 10137
rect 26000 10064 26006 10098
rect 25975 10025 26006 10064
rect 26000 9991 26006 10025
rect 25975 9952 26006 9991
rect 26000 9918 26006 9952
rect 25975 9879 26006 9918
rect 26000 9845 26006 9879
rect 25975 9806 26006 9845
rect 1289 9788 1545 9795
rect 1289 9754 1301 9788
rect 1339 9754 1400 9788
rect 1434 9754 1495 9788
rect 1533 9754 1545 9788
rect 1289 9747 1545 9754
rect 26000 9772 26006 9806
rect 1073 9671 1083 9710
rect 25975 9733 26006 9772
rect 893 9599 903 9638
rect 1077 9637 1083 9671
rect 893 9565 899 9599
rect 1073 9598 1083 9637
rect 893 9526 903 9565
rect 1077 9564 1083 9598
rect 893 9492 899 9526
rect 1073 9525 1083 9564
rect 893 9453 903 9492
rect 1077 9491 1083 9525
rect 893 9419 899 9453
rect 1073 9452 1083 9491
rect 893 9380 903 9419
rect 1077 9418 1083 9452
rect 893 9346 899 9380
rect 1073 9379 1083 9418
rect 893 9307 903 9346
rect 1077 9345 1083 9379
rect 893 9273 899 9307
rect 1073 9306 1083 9345
rect 893 9234 903 9273
rect 1077 9272 1083 9306
rect 893 9200 899 9234
rect 1073 9233 1083 9272
rect 893 9161 903 9200
rect 1077 9199 1083 9233
rect 893 9127 899 9161
rect 1073 9160 1083 9199
rect 1244 9691 1278 9703
rect 1244 9619 1278 9653
rect 1244 9551 1278 9584
rect 1244 9483 1278 9510
rect 1244 9415 1278 9449
rect 1244 9347 1278 9381
rect 1244 9279 1278 9313
rect 1244 9211 1278 9245
rect 1244 9161 1278 9177
rect 1400 9687 1434 9703
rect 1400 9619 1434 9653
rect 1400 9551 1434 9585
rect 1400 9483 1434 9517
rect 1400 9415 1434 9420
rect 1400 9347 1434 9348
rect 1400 9279 1434 9313
rect 1400 9211 1434 9245
rect 1400 9161 1434 9177
rect 1556 9691 1590 9703
rect 1556 9619 1590 9653
rect 1556 9551 1590 9584
rect 1556 9483 1590 9510
rect 1556 9415 1590 9449
rect 1556 9347 1590 9381
rect 1556 9279 1590 9313
rect 1556 9211 1590 9245
rect 1556 9161 1590 9177
rect 26000 9699 26006 9733
rect 25975 9660 26006 9699
rect 26000 9626 26006 9660
rect 25975 9587 26006 9626
rect 26000 9553 26006 9587
rect 25975 9514 26006 9553
rect 26000 9480 26006 9514
rect 25975 9441 26006 9480
rect 26000 9407 26006 9441
rect 25975 9368 26006 9407
rect 26000 9334 26006 9368
rect 25975 9295 26006 9334
rect 26000 9261 26006 9295
rect 25975 9222 26006 9261
rect 26000 9188 26006 9222
rect 893 9088 903 9127
rect 1077 9126 1083 9160
rect 893 9054 899 9088
rect 1073 9087 1083 9126
rect 893 9015 903 9054
rect 1077 9053 1083 9087
rect 893 8981 899 9015
rect 1073 9014 1083 9053
rect 893 8942 903 8981
rect 1077 8980 1083 9014
rect 893 8908 899 8942
rect 1073 8941 1083 8980
rect 893 8869 903 8908
rect 1077 8907 1083 8941
rect 893 8835 899 8869
rect 1073 8868 1083 8907
rect 893 8796 903 8835
rect 1077 8834 1083 8868
rect 893 8762 899 8796
rect 1073 8795 1083 8834
rect 893 8723 903 8762
rect 1077 8761 1083 8795
rect 893 8689 899 8723
rect 1073 8722 1083 8761
rect 893 8650 903 8689
rect 1077 8688 1083 8722
rect 893 8616 899 8650
rect 1073 8649 1083 8688
rect 893 8577 903 8616
rect 1077 8615 1083 8649
rect 893 8543 899 8577
rect 1073 8576 1083 8615
rect 893 8504 903 8543
rect 1077 8542 1083 8576
rect 893 8470 899 8504
rect 1073 8503 1083 8542
rect 893 8431 903 8470
rect 1077 8469 1083 8503
rect 893 8397 899 8431
rect 1073 8430 1083 8469
rect 893 8358 903 8397
rect 1077 8396 1083 8430
rect 893 8324 899 8358
rect 1073 8357 1083 8396
rect 893 8285 903 8324
rect 1077 8323 1083 8357
rect 893 8251 899 8285
rect 1073 8284 1083 8323
rect 893 8212 903 8251
rect 1077 8250 1083 8284
rect 893 8178 899 8212
rect 1073 8211 1083 8250
rect 893 8139 903 8178
rect 1077 8177 1083 8211
rect 893 8105 899 8139
rect 1073 8138 1083 8177
rect 25975 9149 26006 9188
rect 26000 9115 26006 9149
rect 25975 9076 26006 9115
rect 26000 9042 26006 9076
rect 25975 9003 26006 9042
rect 26000 8969 26006 9003
rect 25975 8930 26006 8969
rect 26000 8896 26006 8930
rect 25975 8857 26006 8896
rect 26000 8823 26006 8857
rect 25975 8784 26006 8823
rect 26000 8750 26006 8784
rect 25975 8711 26006 8750
rect 26000 8677 26006 8711
rect 25975 8638 26006 8677
rect 26000 8604 26006 8638
rect 25975 8565 26006 8604
rect 26000 8531 26006 8565
rect 25975 8492 26006 8531
rect 26000 8458 26006 8492
rect 25975 8419 26006 8458
rect 26000 8385 26006 8419
rect 25975 8346 26006 8385
rect 26000 8312 26006 8346
rect 25975 8273 26006 8312
rect 26000 8239 26006 8273
rect 25975 8200 26006 8239
rect 893 8066 903 8105
rect 1077 8104 1083 8138
rect 11355 8147 11505 8175
rect 11355 8113 11379 8147
rect 11413 8113 11447 8147
rect 11481 8113 11505 8147
rect 26000 8166 26006 8200
rect 25975 8127 26006 8166
rect 893 8032 899 8066
rect 1073 8065 1083 8104
rect 893 7993 903 8032
rect 1077 8031 1083 8065
rect 893 7959 899 7993
rect 1073 7992 1083 8031
rect 893 7920 903 7959
rect 1077 7958 1083 7992
rect 893 7886 899 7920
rect 1073 7919 1083 7958
rect 893 7847 903 7886
rect 1077 7885 1083 7919
rect 893 7813 899 7847
rect 1073 7846 1083 7885
rect 893 7774 903 7813
rect 1077 7812 1083 7846
rect 893 7740 899 7774
rect 1073 7773 1083 7812
rect 893 7701 903 7740
rect 1077 7739 1083 7773
rect 893 7667 899 7701
rect 1073 7700 1083 7739
rect 893 7628 903 7667
rect 1077 7666 1083 7700
rect 893 7594 899 7628
rect 1073 7627 1083 7666
rect 893 7555 903 7594
rect 1077 7593 1083 7627
rect 893 7521 899 7555
rect 1073 7554 1083 7593
rect 893 7482 903 7521
rect 1077 7520 1083 7554
rect 893 7448 899 7482
rect 1073 7481 1083 7520
rect 893 7409 903 7448
rect 1077 7447 1083 7481
rect 893 7375 899 7409
rect 1073 7408 1083 7447
rect 893 7336 903 7375
rect 1077 7374 1083 7408
rect 893 7302 899 7336
rect 1073 7335 1083 7374
rect 893 7295 903 7302
rect 1077 7301 1083 7335
rect 1073 7295 1083 7301
rect 893 7263 1083 7295
rect 893 7229 899 7263
rect 933 7229 971 7263
rect 1005 7262 1083 7263
rect 1005 7229 1043 7262
rect 893 7228 1043 7229
rect 1077 7228 1083 7262
rect 893 7190 1083 7228
rect 893 7156 899 7190
rect 933 7169 971 7190
rect 1005 7189 1083 7190
rect 1005 7169 1043 7189
rect 893 7117 903 7156
rect 1077 7155 1083 7189
rect 893 7083 899 7117
rect 1073 7116 1083 7155
rect 893 7044 903 7083
rect 1077 7082 1083 7116
rect 893 7010 899 7044
rect 1073 7043 1083 7082
rect 893 6971 903 7010
rect 1077 7009 1083 7043
rect 893 6937 899 6971
rect 1073 6970 1083 7009
rect 893 6898 903 6937
rect 1077 6936 1083 6970
rect 893 6864 899 6898
rect 1073 6897 1083 6936
rect 893 6825 903 6864
rect 1077 6863 1083 6897
rect 1005 6830 1083 6863
rect 26000 8093 26006 8127
rect 25975 8054 26006 8093
rect 26000 8020 26006 8054
rect 25975 7981 26006 8020
rect 26000 7947 26006 7981
rect 25975 7908 26006 7947
rect 26000 7874 26006 7908
rect 25975 7835 26006 7874
rect 26000 7801 26006 7835
rect 25975 7762 26006 7801
rect 26000 7728 26006 7762
rect 25975 7689 26006 7728
rect 26000 7655 26006 7689
rect 25975 7616 26006 7655
rect 893 6791 899 6825
rect 1005 6824 25805 6830
rect 1005 6820 1043 6824
rect 25053 6820 25092 6824
rect 25126 6820 25165 6824
rect 25199 6820 25238 6824
rect 25272 6820 25311 6824
rect 25345 6820 25384 6824
rect 25418 6820 25457 6824
rect 25491 6820 25530 6824
rect 25564 6820 25603 6824
rect 25637 6820 25676 6824
rect 25710 6820 25749 6824
rect 933 6791 971 6795
rect 1005 6791 1039 6820
rect 893 6761 1039 6791
rect 893 6752 903 6761
rect 937 6752 1039 6761
rect 25783 6790 25805 6824
rect 25757 6786 25805 6790
rect 25757 6752 25873 6786
rect 893 6718 899 6752
rect 937 6727 971 6752
rect 933 6718 971 6727
rect 893 6646 971 6718
rect 25855 6718 25873 6752
rect 26000 6718 26006 7616
rect 25825 6684 26006 6718
rect 25825 6680 25859 6684
rect 25855 6650 25859 6680
rect 25893 6680 26006 6684
rect 25893 6650 25894 6680
rect 25125 6646 25164 6650
rect 25198 6646 25237 6650
rect 25271 6646 25310 6650
rect 25344 6646 25383 6650
rect 25417 6646 25456 6650
rect 25490 6646 25529 6650
rect 25563 6646 25602 6650
rect 25636 6646 25675 6650
rect 25709 6646 25748 6650
rect 25782 6646 25821 6650
rect 25855 6646 25894 6650
rect 25928 6646 26006 6680
rect 893 6640 26006 6646
rect 26214 12826 26220 12860
rect 26394 12858 26404 12898
rect 26214 12786 26224 12826
rect 26398 12824 26404 12858
rect 26214 12752 26220 12786
rect 26394 12784 26404 12824
rect 26214 12712 26224 12752
rect 26398 12750 26404 12784
rect 26214 12678 26220 12712
rect 26394 12711 26404 12750
rect 26214 12638 26224 12678
rect 26398 12677 26404 12711
rect 26394 12638 26404 12677
rect 26214 12604 26220 12638
rect 26398 12604 26404 12638
rect 26214 12528 26224 12604
rect 26394 12528 26404 12604
rect 26214 12494 26220 12528
rect 26398 12494 26404 12528
rect 26214 12455 26224 12494
rect 26394 12455 26404 12494
rect 26214 12421 26220 12455
rect 26398 12421 26404 12455
rect 26214 12382 26224 12421
rect 26394 12382 26404 12421
rect 26214 12348 26220 12382
rect 26398 12348 26404 12382
rect 26214 12309 26224 12348
rect 26394 12309 26404 12348
rect 26214 12275 26220 12309
rect 26398 12275 26404 12309
rect 26214 12236 26224 12275
rect 26394 12236 26404 12275
rect 26214 12202 26220 12236
rect 26398 12202 26404 12236
rect 26214 12163 26224 12202
rect 26394 12163 26404 12202
rect 507 6558 517 6597
rect 691 6596 697 6630
rect 507 6524 513 6558
rect 687 6557 697 6596
rect 507 6485 517 6524
rect 691 6523 697 6557
rect 507 6451 513 6485
rect 687 6484 697 6523
rect 507 6412 517 6451
rect 691 6450 697 6484
rect 507 6378 513 6412
rect 687 6411 697 6450
rect 507 6339 517 6378
rect 691 6377 697 6411
rect 507 6305 513 6339
rect 687 6338 697 6377
rect 507 6266 517 6305
rect 691 6304 697 6338
rect 507 6232 513 6266
rect 687 6265 697 6304
rect 507 6193 517 6232
rect 691 6231 697 6265
rect 507 6159 513 6193
rect 687 6192 697 6231
rect 507 6120 517 6159
rect 691 6158 697 6192
rect 507 6086 513 6120
rect 687 6119 697 6158
rect 507 6047 517 6086
rect 691 6085 697 6119
rect 507 6013 513 6047
rect 687 6046 697 6085
rect 507 5974 517 6013
rect 691 6012 697 6046
rect 507 5940 513 5974
rect 687 5973 697 6012
rect 507 5901 517 5940
rect 691 5939 697 5973
rect 507 5867 513 5901
rect 687 5900 697 5939
rect 507 5828 517 5867
rect 691 5866 697 5900
rect 687 5851 697 5866
rect 26214 5851 26220 12163
rect 507 5794 513 5828
rect 687 5827 722 5851
rect 756 5827 791 5851
rect 825 5827 860 5851
rect 507 5755 517 5794
rect 619 5783 657 5817
rect 26258 5783 26292 5793
rect 619 5755 654 5783
rect 507 5721 513 5755
rect 547 5721 585 5749
rect 507 5649 585 5721
rect 26398 5721 26404 12163
rect 26107 5649 26146 5681
rect 26180 5649 26219 5681
rect 26253 5649 26292 5681
rect 26326 5649 26404 5721
rect 507 5643 26404 5649
rect 307 5323 342 5357
rect 376 5323 411 5357
rect 445 5323 480 5357
rect 514 5323 549 5357
rect 583 5323 618 5357
rect 652 5323 687 5357
rect 721 5323 756 5357
rect 790 5323 825 5357
rect 859 5323 894 5357
rect 928 5323 963 5357
rect 997 5323 1032 5357
rect 1066 5323 1101 5357
rect 1135 5323 1170 5357
rect 1204 5323 1239 5357
rect 1273 5323 1308 5357
rect 1342 5323 1377 5357
rect 1411 5323 1446 5357
rect 1480 5323 1515 5357
rect 1549 5323 1584 5357
rect 1618 5323 1653 5357
rect 1687 5323 1722 5357
rect 1756 5323 1791 5357
rect 1825 5323 1860 5357
rect 1894 5323 1929 5357
rect 1963 5323 1998 5357
rect 2032 5323 2067 5357
rect 2101 5323 2136 5357
rect 2170 5323 2205 5357
rect 2239 5323 2274 5357
rect 2308 5323 2343 5357
rect 2377 5323 2412 5357
rect 2446 5323 2481 5357
rect 2515 5323 2550 5357
rect 2584 5323 2619 5357
rect 2653 5323 2688 5357
rect 2722 5323 2757 5357
rect 2791 5323 2826 5357
rect 2860 5323 2895 5357
rect 307 5289 2895 5323
rect 69 5255 273 5261
rect 307 5255 342 5289
rect 376 5255 411 5289
rect 445 5255 480 5289
rect 514 5255 549 5289
rect 583 5255 618 5289
rect 652 5255 687 5289
rect 721 5255 756 5289
rect 790 5255 825 5289
rect 859 5255 894 5289
rect 928 5255 963 5289
rect 997 5255 1032 5289
rect 1066 5255 1101 5289
rect 1135 5255 1170 5289
rect 1204 5255 1239 5289
rect 1273 5255 1308 5289
rect 1342 5255 1377 5289
rect 1411 5255 1446 5289
rect 1480 5255 1515 5289
rect 1549 5255 1584 5289
rect 1618 5255 1653 5289
rect 1687 5255 1722 5289
rect 1756 5255 1791 5289
rect 1825 5255 1860 5289
rect 1894 5255 1929 5289
rect 1963 5255 1998 5289
rect 2032 5255 2067 5289
rect 2101 5255 2136 5289
rect 2170 5255 2205 5289
rect 2239 5255 2274 5289
rect 2308 5255 2343 5289
rect 2377 5255 2412 5289
rect 2446 5255 2481 5289
rect 2515 5255 2550 5289
rect 2584 5255 2619 5289
rect 2653 5255 2688 5289
rect 2722 5255 2757 5289
rect 2791 5255 2826 5289
rect 2860 5255 2895 5289
rect 69 5221 2895 5255
rect 69 5187 273 5221
rect 307 5187 342 5221
rect 376 5187 411 5221
rect 445 5187 480 5221
rect 514 5187 549 5221
rect 583 5187 618 5221
rect 652 5187 687 5221
rect 721 5187 756 5221
rect 790 5187 825 5221
rect 859 5187 894 5221
rect 928 5187 963 5221
rect 997 5187 1032 5221
rect 1066 5187 1101 5221
rect 1135 5187 1170 5221
rect 1204 5187 1239 5221
rect 1273 5187 1308 5221
rect 1342 5187 1377 5221
rect 1411 5187 1446 5221
rect 1480 5187 1515 5221
rect 1549 5187 1584 5221
rect 1618 5187 1653 5221
rect 1687 5187 1722 5221
rect 1756 5187 1791 5221
rect 1825 5187 1860 5221
rect 1894 5187 1929 5221
rect 1963 5187 1998 5221
rect 2032 5187 2067 5221
rect 2101 5187 2136 5221
rect 2170 5187 2205 5221
rect 2239 5187 2274 5221
rect 2308 5187 2343 5221
rect 2377 5187 2412 5221
rect 2446 5187 2481 5221
rect 2515 5187 2550 5221
rect 2584 5187 2619 5221
rect 2653 5187 2688 5221
rect 2722 5187 2757 5221
rect 2791 5187 2826 5221
rect 2860 5187 2895 5221
rect 26593 5187 26797 5221
rect 24637 3326 25041 3622
rect -585 3032 -533 3066
rect -499 3032 -447 3066
rect -413 3032 -362 3066
rect -328 3032 -277 3066
rect -619 2988 -243 3032
rect -585 2954 -533 2988
rect -499 2954 -447 2988
rect -413 2954 -362 2988
rect -328 2954 -277 2988
rect -105 3032 -53 3066
rect -19 3032 33 3066
rect 67 3032 118 3066
rect 152 3032 203 3066
rect -139 2988 237 3032
rect -105 2954 -53 2988
rect -19 2954 33 2988
rect 67 2954 118 2988
rect 152 2954 203 2988
rect 380 3032 432 3066
rect 466 3032 518 3066
rect 552 3032 603 3066
rect 637 3032 688 3066
rect 346 2988 722 3032
rect 380 2954 432 2988
rect 466 2954 518 2988
rect 552 2954 603 2988
rect 637 2954 688 2988
rect 24341 3017 24375 3033
rect 24341 2949 24375 2983
rect -1144 2926 -740 2938
rect -1144 2892 -1123 2926
rect -1089 2892 -1035 2926
rect -1001 2892 -948 2926
rect -914 2892 -861 2926
rect -827 2892 -774 2926
rect 24341 2899 24375 2915
rect 24517 2949 24551 2983
rect -1144 2840 -740 2892
rect -1144 2806 -1123 2840
rect -1089 2806 -1035 2840
rect -1001 2806 -948 2840
rect -914 2806 -861 2840
rect -827 2806 -774 2840
rect -1144 2802 -740 2806
rect 24039 2825 24680 2842
rect 24039 2791 24406 2825
rect 24440 2791 24480 2825
rect 24514 2791 24554 2825
rect 24588 2791 24628 2825
rect 24662 2791 24680 2825
rect 24039 2776 24680 2791
rect 6507 2705 6541 2721
rect 6507 2655 6541 2671
rect 6763 2705 6797 2721
rect 6763 2655 6797 2671
rect 24341 2699 24375 2715
rect 24341 2631 24375 2665
rect 24341 2563 24375 2597
rect 24341 2513 24375 2529
rect 24517 2643 24551 2665
rect 24517 2563 24551 2597
rect 24517 2513 24551 2529
rect 24693 2699 24727 2715
rect 24693 2631 24727 2665
rect 24693 2563 24727 2597
rect 24693 2513 24727 2529
rect -1144 1294 749 1464
rect -1144 1260 -1132 1294
rect -1098 1260 -1058 1294
rect -1024 1260 -984 1294
rect -950 1260 -910 1294
rect -876 1260 -836 1294
rect -802 1260 -762 1294
rect -728 1260 -688 1294
rect -654 1260 -614 1294
rect -580 1260 -540 1294
rect -506 1260 -466 1294
rect -432 1260 -392 1294
rect -358 1260 -319 1294
rect -285 1260 -246 1294
rect -212 1260 -173 1294
rect -139 1260 -100 1294
rect -66 1260 -27 1294
rect 7 1260 46 1294
rect 80 1260 119 1294
rect 153 1260 192 1294
rect 226 1260 265 1294
rect 299 1260 338 1294
rect 372 1260 411 1294
rect 445 1260 484 1294
rect 518 1260 557 1294
rect 591 1260 630 1294
rect 664 1260 703 1294
rect 737 1260 749 1294
rect -1144 1220 749 1260
rect -1144 1186 -1132 1220
rect -1098 1186 -1058 1220
rect -1024 1186 -984 1220
rect -950 1186 -910 1220
rect -876 1186 -836 1220
rect -802 1186 -762 1220
rect -728 1186 -688 1220
rect -654 1186 -614 1220
rect -580 1186 -540 1220
rect -506 1186 -466 1220
rect -432 1186 -392 1220
rect -358 1186 -319 1220
rect -285 1186 -246 1220
rect -212 1186 -173 1220
rect -139 1186 -100 1220
rect -66 1186 -27 1220
rect 7 1186 46 1220
rect 80 1186 119 1220
rect 153 1186 192 1220
rect 226 1186 265 1220
rect 299 1186 338 1220
rect 372 1186 411 1220
rect 445 1186 484 1220
rect 518 1186 557 1220
rect 591 1186 630 1220
rect 664 1186 703 1220
rect 737 1186 749 1220
rect -1144 1146 749 1186
rect -1144 1112 -1132 1146
rect -1098 1112 -1058 1146
rect -1024 1112 -984 1146
rect -950 1112 -910 1146
rect -876 1112 -836 1146
rect -802 1112 -762 1146
rect -728 1112 -688 1146
rect -654 1112 -614 1146
rect -580 1112 -540 1146
rect -506 1112 -466 1146
rect -432 1112 -392 1146
rect -358 1112 -319 1146
rect -285 1112 -246 1146
rect -212 1112 -173 1146
rect -139 1112 -100 1146
rect -66 1112 -27 1146
rect 7 1112 46 1146
rect 80 1112 119 1146
rect 153 1112 192 1146
rect 226 1112 265 1146
rect 299 1112 338 1146
rect 372 1112 411 1146
rect 445 1112 484 1146
rect 518 1112 557 1146
rect 591 1112 630 1146
rect 664 1112 703 1146
rect 737 1112 749 1146
rect -1144 1072 749 1112
rect -1144 1038 -1132 1072
rect -1098 1038 -1058 1072
rect -1024 1038 -984 1072
rect -950 1038 -910 1072
rect -876 1038 -836 1072
rect -802 1038 -762 1072
rect -728 1038 -688 1072
rect -654 1038 -614 1072
rect -580 1038 -540 1072
rect -506 1038 -466 1072
rect -432 1038 -392 1072
rect -358 1038 -319 1072
rect -285 1038 -246 1072
rect -212 1038 -173 1072
rect -139 1038 -100 1072
rect -66 1038 -27 1072
rect 7 1038 46 1072
rect 80 1038 119 1072
rect 153 1038 192 1072
rect 226 1038 265 1072
rect 299 1038 338 1072
rect 372 1038 411 1072
rect 445 1038 484 1072
rect 518 1038 557 1072
rect 591 1038 630 1072
rect 664 1038 703 1072
rect 737 1038 749 1072
rect -1144 998 749 1038
rect -1144 964 -1132 998
rect -1098 964 -1058 998
rect -1024 964 -984 998
rect -950 964 -910 998
rect -876 964 -836 998
rect -802 964 -762 998
rect -728 964 -688 998
rect -654 964 -614 998
rect -580 964 -540 998
rect -506 964 -466 998
rect -432 964 -392 998
rect -358 964 -319 998
rect -285 964 -246 998
rect -212 964 -173 998
rect -139 964 -100 998
rect -66 964 -27 998
rect 7 964 46 998
rect 80 964 119 998
rect 153 964 192 998
rect 226 964 265 998
rect 299 964 338 998
rect 372 964 411 998
rect 445 964 484 998
rect 518 964 557 998
rect 591 964 630 998
rect 664 964 703 998
rect 737 964 749 998
rect -1144 924 749 964
rect -1144 890 -1132 924
rect -1098 890 -1058 924
rect -1024 890 -984 924
rect -950 890 -910 924
rect -876 890 -836 924
rect -802 890 -762 924
rect -728 890 -688 924
rect -654 890 -614 924
rect -580 890 -540 924
rect -506 890 -466 924
rect -432 890 -392 924
rect -358 890 -319 924
rect -285 890 -246 924
rect -212 890 -173 924
rect -139 890 -100 924
rect -66 890 -27 924
rect 7 890 46 924
rect 80 890 119 924
rect 153 890 192 924
rect 226 890 265 924
rect 299 890 338 924
rect 372 890 411 924
rect 445 890 484 924
rect 518 890 557 924
rect 591 890 630 924
rect 664 890 703 924
rect 737 890 749 924
rect -1144 850 749 890
rect -1144 816 -1132 850
rect -1098 816 -1058 850
rect -1024 816 -984 850
rect -950 816 -910 850
rect -876 816 -836 850
rect -802 816 -762 850
rect -728 816 -688 850
rect -654 816 -614 850
rect -580 816 -540 850
rect -506 816 -466 850
rect -432 816 -392 850
rect -358 816 -319 850
rect -285 816 -246 850
rect -212 816 -173 850
rect -139 816 -100 850
rect -66 816 -27 850
rect 7 816 46 850
rect 80 816 119 850
rect 153 816 192 850
rect 226 816 265 850
rect 299 816 338 850
rect 372 816 411 850
rect 445 816 484 850
rect 518 816 557 850
rect 591 816 630 850
rect 664 816 703 850
rect 737 816 749 850
rect -1144 808 749 816
rect 23701 1193 25860 1199
rect 23701 1159 23779 1193
rect 23814 1159 23848 1193
rect 23886 1159 23916 1193
rect 23959 1159 23984 1193
rect 24032 1159 24052 1193
rect 24105 1159 24120 1193
rect 24178 1159 24188 1193
rect 24251 1159 24256 1193
rect 24358 1159 24363 1193
rect 24426 1159 24436 1193
rect 24494 1159 24509 1193
rect 24562 1159 24582 1193
rect 24630 1159 24655 1193
rect 24698 1159 24728 1193
rect 24766 1159 24800 1193
rect 24835 1159 24868 1193
rect 24908 1159 24936 1193
rect 24981 1159 25004 1193
rect 25054 1159 25072 1193
rect 25127 1159 25140 1193
rect 25200 1159 25208 1193
rect 25273 1159 25276 1193
rect 25310 1159 25312 1193
rect 25378 1159 25385 1193
rect 25446 1159 25458 1193
rect 25514 1159 25531 1193
rect 25582 1159 25604 1193
rect 25650 1159 25676 1193
rect 25718 1159 25748 1193
rect 25786 1159 25860 1193
rect 23701 1153 25860 1159
rect 23701 1125 23747 1153
rect 23701 1071 23707 1125
rect 23741 1071 23747 1125
rect 25814 1125 25860 1153
rect 23701 1057 23747 1071
rect 23701 1023 23707 1057
rect 23741 1023 23747 1057
rect 24460 1076 24500 1110
rect 24534 1076 24574 1110
rect 24608 1076 24648 1110
rect 24164 1027 24229 1029
rect 24263 1027 24328 1029
rect 24426 1027 24682 1076
rect 25220 1076 25260 1110
rect 25294 1076 25334 1110
rect 25368 1076 25408 1110
rect 24933 1027 24992 1029
rect 25026 1027 25084 1029
rect 25186 1027 25442 1076
rect 23701 989 23747 1023
rect 24114 993 24130 1027
rect 24164 993 24225 1027
rect 24263 995 24320 1027
rect 24362 995 24370 1027
rect 24259 993 24320 995
rect 24354 993 24370 995
rect 24426 993 24442 1027
rect 24476 993 24537 1027
rect 24571 993 24632 1027
rect 24666 993 24682 1027
rect 24874 993 24890 1027
rect 24933 995 24985 1027
rect 25026 995 25080 1027
rect 25118 995 25130 1027
rect 24924 993 24985 995
rect 25019 993 25080 995
rect 25114 993 25130 995
rect 25186 993 25202 1027
rect 25236 993 25297 1027
rect 25331 993 25392 1027
rect 25426 993 25442 1027
rect 25814 1087 25820 1125
rect 25854 1087 25860 1125
rect 25814 1057 25860 1087
rect 25814 1008 25820 1057
rect 25854 1008 25860 1057
rect 23701 945 23707 989
rect 23741 945 23747 989
rect 25814 989 25860 1008
rect 23701 921 23747 945
rect 23701 859 23707 921
rect 23741 859 23747 921
rect 23701 853 23747 859
rect 23701 819 23707 853
rect 23741 819 23747 853
rect 24069 934 24103 949
rect 24225 948 24259 949
rect 24090 933 24128 934
rect 24103 900 24128 933
rect 24215 933 24279 948
rect 24381 934 24415 949
rect 23953 873 23987 885
rect 24069 883 24103 899
rect 24215 899 24225 933
rect 24259 899 24279 933
rect 24381 933 24419 934
rect 23701 807 23747 819
rect 23701 751 23707 807
rect 23741 751 23747 807
rect 24215 836 24279 899
rect 24415 900 24419 933
rect 24522 933 24586 949
rect 24693 934 24727 949
rect 24381 883 24415 899
rect 24522 899 24537 933
rect 24571 899 24586 933
rect 24664 933 24702 934
rect 24664 900 24693 933
rect 24829 907 24863 923
rect 24522 836 24586 899
rect 24693 883 24727 899
rect 24249 802 24287 836
rect 24511 802 24549 836
rect 24583 802 24586 836
rect 24971 907 25009 927
rect 24971 893 24985 907
rect 25141 907 25175 923
rect 24829 834 24863 872
rect 24985 857 25019 873
rect 25311 907 25349 927
rect 25331 893 25349 907
rect 25453 907 25487 923
rect 25175 873 25179 893
rect 25141 859 25179 873
rect 25141 857 25175 859
rect 25297 857 25331 873
rect 25569 919 25603 938
rect 25569 861 25603 866
rect 25814 929 25820 989
rect 25854 929 25860 989
rect 25814 921 25860 929
rect 25814 887 25820 921
rect 25854 887 25860 921
rect 25814 884 25860 887
rect 25453 818 25487 856
rect 25814 819 25820 884
rect 25854 819 25860 884
rect 25814 805 25860 819
rect 23701 721 23747 751
rect 23701 687 23707 721
rect 23741 687 23747 721
rect 23701 655 23747 687
rect 25814 751 25820 805
rect 25854 751 25860 805
rect 25814 727 25860 751
rect 25814 683 25820 727
rect 25854 683 25860 727
rect 25814 655 25860 683
rect 23701 649 25860 655
rect 23701 615 23775 649
rect 23813 615 23843 649
rect 23885 615 23911 649
rect 23957 615 23979 649
rect 24030 615 24047 649
rect 24103 615 24115 649
rect 24176 615 24183 649
rect 24249 615 24251 649
rect 24285 615 24288 649
rect 24353 615 24361 649
rect 24421 615 24434 649
rect 24489 615 24507 649
rect 24557 615 24580 649
rect 24625 615 24653 649
rect 24693 615 24726 649
rect 24761 615 24795 649
rect 24833 615 24863 649
rect 24906 615 24931 649
rect 24979 615 24999 649
rect 25052 615 25067 649
rect 25125 615 25135 649
rect 25198 615 25203 649
rect 25305 615 25310 649
rect 25373 615 25383 649
rect 25441 615 25456 649
rect 25509 615 25529 649
rect 25577 615 25602 649
rect 25645 615 25675 649
rect 25713 615 25747 649
rect 25782 615 25860 649
rect 23701 609 25860 615
<< viali >>
rect 1174 22665 1208 22667
rect 1174 22633 1208 22665
rect 1252 22633 1286 22667
rect 1330 22665 1364 22667
rect 1408 22665 1442 22667
rect 1486 22665 1520 22667
rect 1564 22665 1598 22667
rect 1642 22665 1676 22667
rect 1720 22665 1754 22667
rect 1330 22633 1364 22665
rect 1408 22633 1442 22665
rect 1486 22633 1520 22665
rect 1564 22633 1598 22665
rect 1642 22633 1676 22665
rect 1720 22633 1754 22665
rect 1096 22561 1098 22595
rect 1098 22561 1130 22595
rect 1168 22561 1200 22595
rect 1200 22561 1202 22595
rect 1252 22561 1286 22595
rect 1330 22563 1364 22595
rect 1408 22563 1442 22595
rect 1486 22563 1520 22595
rect 1564 22563 1598 22595
rect 1642 22563 1676 22595
rect 1720 22563 1756 22595
rect 1756 22584 1826 22595
rect 1756 22563 1790 22584
rect 1330 22561 1364 22563
rect 1408 22561 1442 22563
rect 1486 22561 1520 22563
rect 1564 22561 1598 22563
rect 1642 22561 1676 22563
rect 1096 22488 1098 22522
rect 1098 22488 1130 22522
rect 1168 22488 1200 22522
rect 1200 22488 1202 22522
rect 1096 22415 1098 22449
rect 1098 22415 1130 22449
rect 1168 22415 1200 22449
rect 1200 22415 1202 22449
rect 1720 22550 1790 22563
rect 1790 22550 1824 22584
rect 1824 22550 1826 22584
rect 1720 22516 1826 22550
rect 1720 22489 1722 22516
rect 1722 22489 1824 22516
rect 1824 22489 1826 22516
rect 1720 22416 1722 22450
rect 1722 22416 1754 22450
rect 1792 22416 1824 22450
rect 1824 22416 1826 22450
rect 1096 22342 1098 22376
rect 1098 22342 1130 22376
rect 1168 22342 1200 22376
rect 1200 22342 1202 22376
rect 1366 22370 1400 22393
rect 1096 22269 1098 22303
rect 1098 22269 1130 22303
rect 1168 22269 1200 22303
rect 1200 22269 1202 22303
rect 1366 22359 1400 22370
rect 1522 22370 1556 22393
rect 1366 22287 1400 22321
rect 1522 22359 1556 22370
rect 1522 22287 1556 22321
rect 1720 22343 1722 22377
rect 1722 22343 1754 22377
rect 1792 22343 1824 22377
rect 1824 22343 1826 22377
rect 1720 22270 1722 22304
rect 1722 22270 1754 22304
rect 1792 22270 1824 22304
rect 1824 22270 1826 22304
rect 1096 22196 1098 22230
rect 1098 22196 1130 22230
rect 1168 22196 1200 22230
rect 1200 22196 1202 22230
rect 1096 22123 1098 22157
rect 1098 22123 1130 22157
rect 1168 22123 1200 22157
rect 1200 22123 1202 22157
rect 1096 22050 1098 22084
rect 1098 22050 1130 22084
rect 1168 22050 1200 22084
rect 1200 22050 1202 22084
rect 1096 21977 1098 22011
rect 1098 21977 1130 22011
rect 1168 21977 1200 22011
rect 1200 21977 1202 22011
rect 1096 16783 1098 21938
rect 1098 16783 1200 21938
rect 1200 16783 1202 21938
rect 1096 16749 1202 16783
rect 1096 16511 1098 16749
rect 1098 16511 1200 16749
rect 1200 16511 1202 16749
rect 1096 16477 1202 16511
rect 1096 16443 1098 16477
rect 1098 16443 1132 16477
rect 1132 16464 1202 16477
rect 1288 22243 1322 22255
rect 1288 22221 1322 22243
rect 1288 22175 1322 22183
rect 1288 22149 1322 22175
rect 1288 22107 1322 22111
rect 1288 22077 1322 22107
rect 1288 22005 1322 22039
rect 1288 21937 1322 21967
rect 1288 21933 1322 21937
rect 1288 21869 1322 21895
rect 1288 21861 1322 21869
rect 1288 21801 1322 21823
rect 1288 21789 1322 21801
rect 1288 21733 1322 21751
rect 1288 21717 1322 21733
rect 1444 22243 1478 22255
rect 1444 22221 1478 22243
rect 1444 22175 1478 22183
rect 1444 22149 1478 22175
rect 1444 22107 1478 22111
rect 1444 22077 1478 22107
rect 1444 22005 1478 22039
rect 1444 21937 1478 21967
rect 1444 21933 1478 21937
rect 1444 21869 1478 21895
rect 1444 21861 1478 21869
rect 1444 21801 1478 21823
rect 1444 21789 1478 21801
rect 1444 21733 1478 21751
rect 1444 21717 1478 21733
rect 1600 22243 1634 22255
rect 1600 22221 1634 22243
rect 1600 22175 1634 22183
rect 1600 22149 1634 22175
rect 1600 22107 1634 22111
rect 1600 22077 1634 22107
rect 1600 22005 1634 22039
rect 1600 21937 1634 21967
rect 1600 21933 1634 21937
rect 1600 21869 1634 21895
rect 1600 21861 1634 21869
rect 1600 21801 1634 21823
rect 1600 21789 1634 21801
rect 1600 21733 1634 21751
rect 1600 21717 1634 21733
rect 1720 22197 1722 22231
rect 1722 22197 1754 22231
rect 1792 22197 1824 22231
rect 1824 22197 1826 22231
rect 1720 22124 1722 22158
rect 1722 22124 1754 22158
rect 1792 22124 1824 22158
rect 1824 22124 1826 22158
rect 1720 22051 1722 22085
rect 1722 22051 1754 22085
rect 1792 22051 1824 22085
rect 1824 22051 1826 22085
rect 1720 21978 1722 22012
rect 1722 21978 1754 22012
rect 1792 21978 1824 22012
rect 1824 21978 1826 22012
rect 1720 21905 1722 21939
rect 1722 21905 1754 21939
rect 1792 21905 1824 21939
rect 1824 21905 1826 21939
rect 1720 21832 1722 21866
rect 1722 21832 1754 21866
rect 1792 21832 1824 21866
rect 1824 21832 1826 21866
rect 1720 21759 1722 21793
rect 1722 21759 1754 21793
rect 1792 21759 1824 21793
rect 1824 21759 1826 21793
rect 1366 21674 1400 21708
rect 1366 21602 1400 21636
rect 1522 21674 1556 21708
rect 1720 21686 1722 21720
rect 1722 21686 1754 21720
rect 1792 21686 1824 21720
rect 1824 21686 1826 21720
rect 1522 21602 1556 21636
rect 1720 21613 1722 21647
rect 1722 21613 1754 21647
rect 1792 21613 1824 21647
rect 1824 21613 1826 21647
rect 1288 21577 1322 21593
rect 1288 21559 1322 21577
rect 1288 21509 1322 21521
rect 1288 21487 1322 21509
rect 1288 21441 1322 21449
rect 1288 21415 1322 21441
rect 1288 21373 1322 21377
rect 1288 21343 1322 21373
rect 1288 21271 1322 21305
rect 1288 21203 1322 21233
rect 1288 21199 1322 21203
rect 1288 21135 1322 21161
rect 1288 21127 1322 21135
rect 1288 21067 1322 21089
rect 1288 21055 1322 21067
rect 1444 21577 1478 21593
rect 1444 21559 1478 21577
rect 1444 21509 1478 21521
rect 1444 21487 1478 21509
rect 1444 21441 1478 21449
rect 1444 21415 1478 21441
rect 1444 21373 1478 21377
rect 1444 21343 1478 21373
rect 1444 21271 1478 21305
rect 1444 21203 1478 21233
rect 1444 21199 1478 21203
rect 1444 21135 1478 21161
rect 1444 21127 1478 21135
rect 1444 21067 1478 21089
rect 1444 21055 1478 21067
rect 1600 21577 1634 21593
rect 1600 21559 1634 21577
rect 1600 21509 1634 21521
rect 1600 21487 1634 21509
rect 1600 21441 1634 21449
rect 1600 21415 1634 21441
rect 1600 21373 1634 21377
rect 1600 21343 1634 21373
rect 1600 21271 1634 21305
rect 1600 21203 1634 21233
rect 1600 21199 1634 21203
rect 1600 21135 1634 21161
rect 1600 21127 1634 21135
rect 1600 21067 1634 21089
rect 1720 21540 1722 21574
rect 1722 21540 1754 21574
rect 1792 21540 1824 21574
rect 1824 21540 1826 21574
rect 1720 21467 1722 21501
rect 1722 21467 1754 21501
rect 1792 21467 1824 21501
rect 1824 21467 1826 21501
rect 1720 21394 1722 21428
rect 1722 21394 1754 21428
rect 1792 21394 1824 21428
rect 1824 21394 1826 21428
rect 1720 21321 1722 21355
rect 1722 21321 1754 21355
rect 1792 21321 1824 21355
rect 1824 21321 1826 21355
rect 1720 21248 1722 21282
rect 1722 21248 1754 21282
rect 1792 21248 1824 21282
rect 1824 21248 1826 21282
rect 1720 21175 1722 21209
rect 1722 21175 1754 21209
rect 1792 21175 1824 21209
rect 1824 21175 1826 21209
rect 1720 21102 1722 21136
rect 1722 21102 1754 21136
rect 1792 21102 1824 21136
rect 1824 21102 1826 21136
rect 1600 21055 1634 21067
rect 1244 16464 1278 16466
rect 1320 16464 1354 16466
rect 1395 16464 1429 16466
rect 1470 16464 1504 16466
rect 1545 16464 1579 16466
rect 1620 16464 1654 16466
rect 1132 16443 1166 16464
rect 1096 16432 1166 16443
rect 1166 16432 1202 16464
rect 1244 16432 1278 16464
rect 1320 16432 1354 16464
rect 1395 16432 1429 16464
rect 1470 16432 1504 16464
rect 1545 16432 1579 16464
rect 1620 16432 1654 16464
rect 1695 16432 1722 16466
rect 1722 16432 1729 16466
rect 1168 16362 1202 16394
rect 1246 16362 1280 16394
rect 1324 16362 1358 16394
rect 1402 16362 1436 16394
rect 1480 16362 1514 16394
rect 1558 16362 1592 16394
rect 1636 16362 1670 16394
rect 1714 16362 1744 16394
rect 1744 16362 1748 16394
rect 1792 16383 1826 16417
rect 1168 16360 1202 16362
rect 1246 16360 1280 16362
rect 1324 16360 1358 16362
rect 1402 16360 1436 16362
rect 1480 16360 1514 16362
rect 1558 16360 1592 16362
rect 1636 16360 1670 16362
rect 1714 16360 1748 16362
rect 585 13222 619 13226
rect 658 13222 692 13226
rect 731 13222 765 13226
rect 804 13222 26326 13226
rect 585 13192 619 13222
rect 658 13192 692 13222
rect 731 13192 765 13222
rect 513 13120 517 13154
rect 517 13120 551 13154
rect 551 13120 585 13154
rect 585 13120 619 13154
rect 658 13120 692 13154
rect 731 13120 765 13154
rect 804 13120 26119 13222
rect 26119 13188 26154 13222
rect 26154 13188 26188 13222
rect 26188 13188 26223 13222
rect 26223 13188 26257 13222
rect 26257 13188 26292 13222
rect 26292 13188 26326 13222
rect 26119 13154 26326 13188
rect 26119 13120 26154 13154
rect 26154 13120 26188 13154
rect 26188 13120 26223 13154
rect 26223 13120 26257 13154
rect 26257 13120 26292 13154
rect 26292 13120 26326 13154
rect 26364 13120 26394 13154
rect 26394 13120 26398 13154
rect 513 13085 619 13120
rect 513 13051 517 13085
rect 517 13051 551 13085
rect 551 13051 585 13085
rect 585 13051 619 13085
rect 619 13052 653 13082
rect 653 13052 691 13082
rect 730 13052 764 13082
rect 803 13052 837 13082
rect 876 13052 26051 13120
rect 26051 13086 26254 13120
rect 26051 13052 26086 13086
rect 26086 13052 26120 13086
rect 26120 13052 26155 13086
rect 26155 13052 26189 13086
rect 26189 13052 26224 13086
rect 619 13051 691 13052
rect 513 13017 691 13051
rect 730 13048 764 13052
rect 803 13048 837 13052
rect 876 13048 26224 13052
rect 26224 13048 26254 13086
rect 26292 13046 26326 13080
rect 26364 13046 26394 13080
rect 26394 13046 26398 13080
rect 513 13016 653 13017
rect 513 12982 517 13016
rect 517 12982 551 13016
rect 551 12982 585 13016
rect 585 12982 619 13016
rect 619 12983 653 13016
rect 653 12983 687 13017
rect 687 12983 691 13017
rect 619 12982 691 12983
rect 513 12948 691 12982
rect 513 12947 653 12948
rect 513 12913 517 12947
rect 517 12913 551 12947
rect 551 12913 585 12947
rect 585 12913 619 12947
rect 619 12914 653 12947
rect 653 12914 687 12948
rect 687 12914 691 12948
rect 619 12913 691 12914
rect 513 12879 691 12913
rect 513 12878 653 12879
rect 513 12844 517 12878
rect 517 12844 551 12878
rect 551 12844 585 12878
rect 585 12844 619 12878
rect 619 12845 653 12878
rect 653 12845 687 12879
rect 687 12845 691 12879
rect 619 12844 691 12845
rect 513 12810 691 12844
rect 513 12809 653 12810
rect 513 12775 517 12809
rect 517 12775 551 12809
rect 551 12775 585 12809
rect 585 12775 619 12809
rect 619 12776 653 12809
rect 653 12776 687 12810
rect 687 12776 691 12810
rect 619 12775 691 12776
rect 513 12741 691 12775
rect 513 12740 653 12741
rect 513 12706 517 12740
rect 517 12706 551 12740
rect 551 12706 585 12740
rect 585 12706 619 12740
rect 619 12707 653 12740
rect 653 12707 687 12741
rect 687 12707 691 12741
rect 619 12706 691 12707
rect 513 12672 691 12706
rect 513 12671 653 12672
rect 513 12637 517 12671
rect 517 12637 551 12671
rect 551 12637 585 12671
rect 585 12637 619 12671
rect 619 12638 653 12671
rect 653 12638 687 12672
rect 687 12638 691 12672
rect 619 12637 691 12638
rect 513 12603 691 12637
rect 513 12602 653 12603
rect 513 12568 517 12602
rect 517 12568 551 12602
rect 551 12568 585 12602
rect 585 12568 619 12602
rect 619 12569 653 12602
rect 653 12569 687 12603
rect 687 12569 691 12603
rect 619 12568 691 12569
rect 513 12534 691 12568
rect 513 12533 653 12534
rect 513 12499 517 12533
rect 517 12499 551 12533
rect 551 12499 585 12533
rect 585 12499 619 12533
rect 619 12500 653 12533
rect 653 12500 687 12534
rect 687 12500 691 12534
rect 619 12499 691 12500
rect 513 12465 691 12499
rect 513 12464 653 12465
rect 513 12430 517 12464
rect 517 12430 551 12464
rect 551 12430 585 12464
rect 585 12430 619 12464
rect 619 12431 653 12464
rect 653 12431 687 12465
rect 687 12431 691 12465
rect 619 12430 691 12431
rect 513 12396 691 12430
rect 513 12395 653 12396
rect 513 12361 517 12395
rect 517 12361 551 12395
rect 551 12361 585 12395
rect 585 12361 619 12395
rect 619 12362 653 12395
rect 653 12362 687 12396
rect 687 12362 691 12396
rect 619 12361 691 12362
rect 513 12327 691 12361
rect 513 12326 653 12327
rect 513 12292 517 12326
rect 517 12292 551 12326
rect 551 12292 585 12326
rect 585 12292 619 12326
rect 619 12293 653 12326
rect 653 12293 687 12327
rect 687 12293 691 12327
rect 619 12292 691 12293
rect 513 12258 691 12292
rect 513 12257 653 12258
rect 513 12223 517 12257
rect 517 12223 551 12257
rect 551 12223 585 12257
rect 585 12223 619 12257
rect 619 12224 653 12257
rect 653 12224 687 12258
rect 687 12224 691 12258
rect 619 12223 691 12224
rect 513 12189 691 12223
rect 513 12188 653 12189
rect 513 12154 517 12188
rect 517 12154 551 12188
rect 551 12154 585 12188
rect 585 12154 619 12188
rect 619 12155 653 12188
rect 653 12155 687 12189
rect 687 12155 691 12189
rect 619 12154 691 12155
rect 513 12120 691 12154
rect 513 12119 653 12120
rect 513 12085 517 12119
rect 517 12085 551 12119
rect 551 12085 585 12119
rect 585 12085 619 12119
rect 619 12086 653 12119
rect 653 12086 687 12120
rect 687 12086 691 12120
rect 619 12085 691 12086
rect 513 12051 691 12085
rect 513 12050 653 12051
rect 513 12016 517 12050
rect 517 12016 551 12050
rect 551 12016 585 12050
rect 585 12016 619 12050
rect 619 12017 653 12050
rect 653 12017 687 12051
rect 687 12017 691 12051
rect 619 12016 691 12017
rect 513 11982 691 12016
rect 513 11981 653 11982
rect 513 11947 517 11981
rect 517 11947 551 11981
rect 551 11947 585 11981
rect 585 11947 619 11981
rect 619 11948 653 11981
rect 653 11948 687 11982
rect 687 11948 691 11982
rect 619 11947 691 11948
rect 513 11913 691 11947
rect 513 11912 653 11913
rect 513 11878 517 11912
rect 517 11878 551 11912
rect 551 11878 585 11912
rect 585 11878 619 11912
rect 619 11879 653 11912
rect 653 11879 687 11913
rect 687 11879 691 11913
rect 619 11878 691 11879
rect 513 11844 691 11878
rect 513 11843 653 11844
rect 513 11809 517 11843
rect 517 11809 551 11843
rect 551 11809 585 11843
rect 585 11809 619 11843
rect 619 11810 653 11843
rect 653 11810 687 11844
rect 687 11810 691 11844
rect 619 11809 691 11810
rect 513 11775 691 11809
rect 513 11774 653 11775
rect 513 11740 517 11774
rect 517 11740 551 11774
rect 551 11740 585 11774
rect 585 11740 619 11774
rect 619 11741 653 11774
rect 653 11741 687 11775
rect 687 11741 691 11775
rect 619 11740 691 11741
rect 513 11706 691 11740
rect 513 11705 653 11706
rect 513 11671 517 11705
rect 517 11671 551 11705
rect 551 11671 585 11705
rect 585 11671 619 11705
rect 619 11672 653 11705
rect 653 11672 687 11706
rect 687 11672 691 11706
rect 619 11671 691 11672
rect 513 11637 691 11671
rect 513 11636 653 11637
rect 513 11602 517 11636
rect 517 11602 551 11636
rect 551 11602 585 11636
rect 585 11602 619 11636
rect 619 11603 653 11636
rect 653 11603 687 11637
rect 687 11603 691 11637
rect 619 11602 691 11603
rect 513 11568 691 11602
rect 513 11567 653 11568
rect 513 11533 517 11567
rect 517 11533 551 11567
rect 551 11533 585 11567
rect 585 11533 619 11567
rect 619 11534 653 11567
rect 653 11534 687 11568
rect 687 11534 691 11568
rect 619 11533 691 11534
rect 513 11499 691 11533
rect 513 11498 653 11499
rect 513 11464 517 11498
rect 517 11464 551 11498
rect 551 11464 585 11498
rect 585 11464 619 11498
rect 619 11465 653 11498
rect 653 11465 687 11499
rect 687 11465 691 11499
rect 619 11464 691 11465
rect 513 11430 691 11464
rect 513 11429 653 11430
rect 513 11395 517 11429
rect 517 11395 551 11429
rect 551 11395 585 11429
rect 585 11395 619 11429
rect 619 11396 653 11429
rect 653 11396 687 11430
rect 687 11396 691 11430
rect 619 11395 691 11396
rect 513 11361 691 11395
rect 513 11360 653 11361
rect 513 11326 517 11360
rect 517 11326 551 11360
rect 551 11326 585 11360
rect 585 11326 619 11360
rect 619 11327 653 11360
rect 653 11327 687 11361
rect 687 11327 691 11361
rect 619 11326 691 11327
rect 513 11292 691 11326
rect 513 11291 653 11292
rect 513 11257 517 11291
rect 517 11257 551 11291
rect 551 11257 585 11291
rect 585 11257 619 11291
rect 619 11258 653 11291
rect 653 11258 687 11292
rect 687 11258 691 11292
rect 619 11257 691 11258
rect 513 11223 691 11257
rect 513 11222 653 11223
rect 513 11188 517 11222
rect 517 11188 551 11222
rect 551 11188 585 11222
rect 585 11188 619 11222
rect 619 11189 653 11222
rect 653 11189 687 11223
rect 687 11189 691 11223
rect 619 11188 691 11189
rect 513 11154 691 11188
rect 513 11153 653 11154
rect 513 11119 517 11153
rect 517 11119 551 11153
rect 551 11119 585 11153
rect 585 11119 619 11153
rect 619 11120 653 11153
rect 653 11120 687 11154
rect 687 11120 691 11154
rect 619 11119 691 11120
rect 513 11085 691 11119
rect 513 11084 653 11085
rect 513 11050 517 11084
rect 517 11050 551 11084
rect 551 11050 585 11084
rect 585 11050 619 11084
rect 619 11051 653 11084
rect 653 11051 687 11085
rect 687 11051 691 11085
rect 619 11050 691 11051
rect 513 11016 691 11050
rect 513 11015 653 11016
rect 513 10981 517 11015
rect 517 10981 551 11015
rect 551 10981 585 11015
rect 585 10981 619 11015
rect 619 10982 653 11015
rect 653 10982 687 11016
rect 687 10982 691 11016
rect 619 10981 691 10982
rect 513 10947 691 10981
rect 513 10946 653 10947
rect 513 10912 517 10946
rect 517 10912 551 10946
rect 551 10912 585 10946
rect 585 10912 619 10946
rect 619 10913 653 10946
rect 653 10913 687 10947
rect 687 10913 691 10947
rect 619 10912 691 10913
rect 513 10878 691 10912
rect 513 10877 653 10878
rect 513 10843 517 10877
rect 517 10843 551 10877
rect 551 10843 585 10877
rect 585 10843 619 10877
rect 619 10844 653 10877
rect 653 10844 687 10878
rect 687 10844 691 10878
rect 619 10843 691 10844
rect 513 10809 691 10843
rect 513 10808 653 10809
rect 513 10774 517 10808
rect 517 10774 551 10808
rect 551 10774 585 10808
rect 585 10774 619 10808
rect 619 10775 653 10808
rect 653 10775 687 10809
rect 687 10775 691 10809
rect 619 10774 691 10775
rect 513 10740 691 10774
rect 513 10739 653 10740
rect 513 10705 517 10739
rect 517 10705 551 10739
rect 551 10705 585 10739
rect 585 10705 619 10739
rect 619 10706 653 10739
rect 653 10706 687 10740
rect 687 10706 691 10740
rect 619 10705 691 10706
rect 513 10671 691 10705
rect 513 10670 653 10671
rect 513 10636 517 10670
rect 517 10636 551 10670
rect 551 10636 585 10670
rect 585 10636 619 10670
rect 619 10637 653 10670
rect 653 10637 687 10671
rect 687 10637 691 10671
rect 619 10636 691 10637
rect 513 10602 691 10636
rect 513 10601 653 10602
rect 513 10567 517 10601
rect 517 10567 551 10601
rect 551 10567 585 10601
rect 585 10567 619 10601
rect 619 10568 653 10601
rect 653 10568 687 10602
rect 687 10568 691 10602
rect 619 10567 691 10568
rect 513 10533 691 10567
rect 513 10532 653 10533
rect 513 10498 517 10532
rect 517 10498 551 10532
rect 551 10498 585 10532
rect 585 10498 619 10532
rect 619 10499 653 10532
rect 653 10499 687 10533
rect 687 10499 691 10533
rect 619 10498 691 10499
rect 513 10464 691 10498
rect 513 10463 653 10464
rect 513 10429 517 10463
rect 517 10429 551 10463
rect 551 10429 585 10463
rect 585 10429 619 10463
rect 619 10430 653 10463
rect 653 10430 687 10464
rect 687 10430 691 10464
rect 619 10429 691 10430
rect 513 10395 691 10429
rect 513 10394 653 10395
rect 513 9816 517 10394
rect 517 10326 619 10394
rect 619 10361 653 10394
rect 653 10361 687 10395
rect 687 10361 691 10395
rect 619 10326 691 10361
rect 517 9816 687 10326
rect 687 9816 691 10326
rect 513 9808 691 9816
rect 26220 12974 26224 13008
rect 26224 12974 26254 13008
rect 26292 12972 26326 13006
rect 26364 12972 26394 13006
rect 26394 12972 26398 13006
rect 26220 12900 26224 12934
rect 26224 12900 26254 12934
rect 26292 12898 26326 12932
rect 26364 12898 26394 12932
rect 26394 12898 26398 12932
rect 513 9748 619 9808
rect 657 9748 691 9769
rect 513 9736 517 9748
rect 517 9736 551 9748
rect 551 9736 585 9748
rect 585 9736 619 9748
rect 657 9735 687 9748
rect 687 9735 691 9748
rect 513 9679 547 9697
rect 585 9679 619 9697
rect 657 9679 691 9696
rect 513 9663 517 9679
rect 517 9663 547 9679
rect 585 9663 619 9679
rect 657 9662 687 9679
rect 687 9662 691 9679
rect 513 9610 547 9624
rect 585 9610 619 9624
rect 657 9610 691 9623
rect 513 9590 517 9610
rect 517 9590 547 9610
rect 585 9590 619 9610
rect 657 9589 687 9610
rect 687 9589 691 9610
rect 513 9541 547 9551
rect 585 9541 619 9551
rect 657 9541 691 9550
rect 513 9517 517 9541
rect 517 9517 547 9541
rect 585 9517 619 9541
rect 657 9516 687 9541
rect 687 9516 691 9541
rect 513 9472 547 9478
rect 585 9472 619 9478
rect 657 9472 691 9477
rect 513 9444 517 9472
rect 517 9444 547 9472
rect 585 9444 619 9472
rect 657 9443 687 9472
rect 687 9443 691 9472
rect 513 9403 547 9405
rect 585 9403 619 9405
rect 657 9403 691 9404
rect 513 9371 517 9403
rect 517 9371 547 9403
rect 585 9371 619 9403
rect 657 9370 687 9403
rect 687 9370 691 9403
rect 513 9300 517 9332
rect 517 9300 547 9332
rect 585 9300 619 9332
rect 657 9300 687 9331
rect 687 9300 691 9331
rect 513 9298 547 9300
rect 585 9298 619 9300
rect 657 9297 691 9300
rect 513 9231 517 9259
rect 517 9231 547 9259
rect 585 9231 619 9259
rect 657 9231 687 9258
rect 687 9231 691 9258
rect 513 9225 547 9231
rect 585 9225 619 9231
rect 657 9224 691 9231
rect 513 9162 517 9186
rect 517 9162 547 9186
rect 585 9162 619 9186
rect 657 9162 687 9185
rect 687 9162 691 9185
rect 513 9152 547 9162
rect 585 9152 619 9162
rect 657 9151 691 9162
rect 513 9093 517 9113
rect 517 9093 547 9113
rect 585 9093 619 9113
rect 657 9093 687 9112
rect 687 9093 691 9112
rect 513 9079 547 9093
rect 585 9079 619 9093
rect 657 9078 691 9093
rect 513 9024 517 9040
rect 517 9024 547 9040
rect 585 9024 619 9040
rect 657 9024 687 9039
rect 687 9024 691 9039
rect 513 9006 547 9024
rect 585 9006 619 9024
rect 657 9005 691 9024
rect 513 8955 517 8967
rect 517 8955 547 8967
rect 585 8955 619 8967
rect 657 8955 687 8966
rect 687 8955 691 8966
rect 513 8933 547 8955
rect 585 8933 619 8955
rect 657 8932 691 8955
rect 513 8886 517 8894
rect 517 8886 547 8894
rect 585 8886 619 8894
rect 657 8886 687 8893
rect 687 8886 691 8893
rect 513 8860 547 8886
rect 585 8860 619 8886
rect 657 8859 691 8886
rect 513 8817 517 8821
rect 517 8817 547 8821
rect 585 8817 619 8821
rect 657 8817 687 8820
rect 687 8817 691 8820
rect 513 8787 547 8817
rect 585 8787 619 8817
rect 657 8786 691 8817
rect 513 8714 547 8748
rect 585 8714 619 8748
rect 657 8713 691 8747
rect 513 8644 547 8675
rect 585 8644 619 8675
rect 657 8644 691 8674
rect 513 8641 517 8644
rect 517 8641 547 8644
rect 585 8641 619 8644
rect 657 8640 687 8644
rect 687 8640 691 8644
rect 513 8575 547 8602
rect 585 8575 619 8602
rect 657 8575 691 8601
rect 513 8568 517 8575
rect 517 8568 547 8575
rect 585 8568 619 8575
rect 657 8567 687 8575
rect 687 8567 691 8575
rect 513 8506 547 8529
rect 585 8506 619 8529
rect 657 8506 691 8528
rect 513 8495 517 8506
rect 517 8495 547 8506
rect 585 8495 619 8506
rect 657 8494 687 8506
rect 687 8494 691 8506
rect 513 8437 547 8456
rect 585 8437 619 8456
rect 657 8437 691 8455
rect 513 8422 517 8437
rect 517 8422 547 8437
rect 585 8422 619 8437
rect 657 8421 687 8437
rect 687 8421 691 8437
rect 513 8368 547 8383
rect 585 8368 619 8383
rect 657 8368 691 8382
rect 513 8349 517 8368
rect 517 8349 547 8368
rect 585 8349 619 8368
rect 657 8348 687 8368
rect 687 8348 691 8368
rect 513 8299 547 8310
rect 585 8299 619 8310
rect 657 8299 691 8309
rect 513 8276 517 8299
rect 517 8276 547 8299
rect 585 8276 619 8299
rect 657 8275 687 8299
rect 687 8275 691 8299
rect 513 8203 517 8237
rect 517 8203 547 8237
rect 585 8203 619 8237
rect 657 8202 687 8236
rect 687 8202 691 8236
rect 513 8130 517 8164
rect 517 8130 547 8164
rect 585 8130 619 8164
rect 657 8129 687 8163
rect 687 8129 691 8163
rect 513 8057 517 8091
rect 517 8057 547 8091
rect 585 8057 619 8091
rect 657 8056 687 8090
rect 687 8056 691 8090
rect 513 7984 517 8018
rect 517 7984 547 8018
rect 585 7984 619 8018
rect 657 7983 687 8017
rect 687 7983 691 8017
rect 513 7911 517 7945
rect 517 7911 547 7945
rect 585 7911 619 7945
rect 657 7910 687 7944
rect 687 7910 691 7944
rect 513 7838 517 7872
rect 517 7838 547 7872
rect 585 7838 619 7872
rect 657 7837 687 7871
rect 687 7837 691 7871
rect 513 7765 517 7799
rect 517 7765 547 7799
rect 585 7765 619 7799
rect 657 7764 687 7798
rect 687 7764 691 7798
rect 513 7692 517 7726
rect 517 7692 547 7726
rect 585 7692 619 7726
rect 657 7691 687 7725
rect 687 7691 691 7725
rect 513 7619 517 7653
rect 517 7619 547 7653
rect 585 7619 619 7653
rect 657 7618 687 7652
rect 687 7618 691 7652
rect 513 7546 517 7580
rect 517 7546 547 7580
rect 585 7546 619 7580
rect 657 7545 687 7579
rect 687 7545 691 7579
rect 513 7473 517 7507
rect 517 7473 547 7507
rect 585 7473 619 7507
rect 657 7472 687 7506
rect 687 7472 691 7506
rect 513 7400 517 7434
rect 517 7400 547 7434
rect 585 7400 619 7434
rect 657 7399 687 7433
rect 687 7399 691 7433
rect 513 7327 517 7361
rect 517 7327 547 7361
rect 585 7327 619 7361
rect 657 7326 687 7360
rect 687 7326 691 7360
rect 513 7254 517 7288
rect 517 7254 547 7288
rect 585 7254 619 7288
rect 657 7253 687 7287
rect 687 7253 691 7287
rect 513 7181 517 7215
rect 517 7181 547 7215
rect 585 7181 619 7215
rect 657 7180 687 7214
rect 687 7180 691 7214
rect 513 7108 517 7142
rect 517 7108 547 7142
rect 585 7108 619 7142
rect 657 7107 687 7141
rect 687 7107 691 7141
rect 513 7035 517 7069
rect 517 7035 547 7069
rect 585 7035 619 7069
rect 657 7034 687 7068
rect 687 7034 691 7068
rect 513 6962 517 6996
rect 517 6962 547 6996
rect 585 6962 619 6996
rect 657 6961 687 6995
rect 687 6961 691 6995
rect 513 6889 517 6923
rect 517 6889 547 6923
rect 585 6889 619 6923
rect 657 6888 687 6922
rect 687 6888 691 6922
rect 513 6816 517 6850
rect 517 6816 547 6850
rect 585 6816 619 6850
rect 657 6815 687 6849
rect 687 6815 691 6849
rect 513 6743 517 6777
rect 517 6743 547 6777
rect 585 6743 619 6777
rect 657 6742 687 6776
rect 687 6742 691 6776
rect 513 6670 517 6704
rect 517 6670 547 6704
rect 585 6670 619 6704
rect 657 6669 687 6703
rect 687 6669 691 6703
rect 513 6597 517 6631
rect 517 6597 547 6631
rect 585 6597 619 6631
rect 971 12837 1005 12840
rect 1044 12837 1078 12840
rect 1117 12837 1151 12840
rect 1190 12837 1224 12840
rect 1263 12837 1297 12840
rect 1336 12837 1370 12840
rect 1409 12837 1443 12840
rect 1482 12837 1516 12840
rect 1555 12837 1589 12840
rect 1628 12837 1662 12840
rect 1701 12837 1735 12840
rect 1774 12837 25928 12840
rect 971 12806 985 12837
rect 985 12806 1005 12837
rect 1044 12806 1053 12837
rect 1053 12806 1078 12837
rect 1117 12806 1151 12837
rect 1190 12806 1224 12837
rect 1263 12806 1297 12837
rect 1336 12806 1370 12837
rect 1409 12806 1443 12837
rect 1482 12806 1516 12837
rect 1555 12806 1589 12837
rect 1628 12806 1662 12837
rect 1701 12806 1735 12837
rect 899 9638 903 12768
rect 903 12696 1005 12768
rect 1044 12735 1053 12768
rect 1053 12735 1078 12768
rect 1117 12735 1151 12768
rect 1044 12734 1078 12735
rect 1117 12734 1121 12735
rect 1121 12734 1151 12735
rect 1190 12734 1224 12768
rect 1263 12734 1297 12768
rect 1336 12734 1370 12768
rect 1409 12734 1443 12768
rect 1482 12734 1516 12768
rect 1555 12734 1589 12768
rect 1628 12734 1662 12768
rect 1701 12734 1735 12768
rect 1774 12735 25907 12837
rect 25907 12735 25928 12837
rect 25966 12736 26000 12768
rect 1774 12734 25839 12735
rect 25839 12734 25928 12735
rect 25966 12734 25975 12736
rect 25975 12734 26000 12736
rect 903 9710 1073 12696
rect 1073 9710 1077 12696
rect 1116 12667 1121 12696
rect 1121 12667 1150 12696
rect 1189 12667 1223 12696
rect 1262 12667 1296 12696
rect 1335 12667 1369 12696
rect 1408 12667 1442 12696
rect 1481 12667 1515 12696
rect 1554 12667 1588 12696
rect 1627 12667 1661 12696
rect 1700 12667 1734 12696
rect 1773 12667 1807 12696
rect 1846 12667 25839 12734
rect 25839 12667 25856 12734
rect 25894 12668 25928 12694
rect 25966 12668 26000 12694
rect 1116 12662 1150 12667
rect 1189 12662 1223 12667
rect 1262 12662 1296 12667
rect 1335 12662 1369 12667
rect 1408 12662 1442 12667
rect 1481 12662 1515 12667
rect 1554 12662 1588 12667
rect 1627 12662 1661 12667
rect 1700 12662 1734 12667
rect 1773 12662 1807 12667
rect 1846 12662 25856 12667
rect 25894 12660 25928 12668
rect 25966 12660 25975 12668
rect 25975 12660 26000 12668
rect 25822 12600 25856 12622
rect 25822 12588 25856 12600
rect 25894 12586 25928 12620
rect 25966 12586 25975 12620
rect 25975 12586 26000 12620
rect 25822 12514 25856 12548
rect 25894 12512 25928 12546
rect 25966 12512 25975 12546
rect 25975 12512 26000 12546
rect 25822 12440 25856 12474
rect 25894 12438 25928 12472
rect 25966 12438 25975 12472
rect 25975 12438 26000 12472
rect 25822 12366 25856 12400
rect 25894 12364 25928 12398
rect 25966 12364 25975 12398
rect 25975 12364 26000 12398
rect 25822 12292 25856 12326
rect 25894 12291 25928 12325
rect 25966 12291 25975 12325
rect 25975 12291 26000 12325
rect 25822 12218 25856 12252
rect 25894 12218 25928 12252
rect 25966 12218 25975 12252
rect 25975 12218 26000 12252
rect 25822 12108 25856 12142
rect 25894 12108 25928 12142
rect 25966 12108 25975 12142
rect 25975 12108 26000 12142
rect 25822 12035 25856 12069
rect 25894 12035 25928 12069
rect 25966 12035 25975 12069
rect 25975 12035 26000 12069
rect 25822 11962 25856 11996
rect 25894 11962 25928 11996
rect 25966 11962 25975 11996
rect 25975 11962 26000 11996
rect 25822 11889 25856 11923
rect 25894 11889 25928 11923
rect 25966 11889 25975 11923
rect 25975 11889 26000 11923
rect 25822 11816 25856 11850
rect 25894 11816 25928 11850
rect 25966 11816 25975 11850
rect 25975 11816 26000 11850
rect 25822 11743 25856 11777
rect 25894 11743 25928 11777
rect 25966 11743 25975 11777
rect 25975 11743 26000 11777
rect 25822 11670 25856 11704
rect 25894 11670 25928 11704
rect 25966 11670 25975 11704
rect 25975 11670 26000 11704
rect 25822 11597 25856 11631
rect 25894 11597 25928 11631
rect 25966 11597 25975 11631
rect 25975 11597 26000 11631
rect 25822 11524 25856 11558
rect 25894 11524 25928 11558
rect 25966 11524 25975 11558
rect 25975 11524 26000 11558
rect 25822 11451 25856 11485
rect 25894 11451 25928 11485
rect 25966 11451 25975 11485
rect 25975 11451 26000 11485
rect 25822 11378 25856 11412
rect 25894 11378 25928 11412
rect 25966 11378 25975 11412
rect 25975 11378 26000 11412
rect 25822 11305 25856 11339
rect 25894 11305 25928 11339
rect 25966 11305 25975 11339
rect 25975 11305 26000 11339
rect 25822 11232 25856 11266
rect 25894 11232 25928 11266
rect 25966 11232 25975 11266
rect 25975 11232 26000 11266
rect 25822 11159 25856 11193
rect 25894 11159 25928 11193
rect 25966 11159 25975 11193
rect 25975 11159 26000 11193
rect 25822 11086 25856 11120
rect 25894 11086 25928 11120
rect 25966 11086 25975 11120
rect 25975 11086 26000 11120
rect 25822 11013 25856 11047
rect 25894 11013 25928 11047
rect 25966 11013 25975 11047
rect 25975 11013 26000 11047
rect 25822 10940 25856 10974
rect 25894 10940 25928 10974
rect 25966 10940 25975 10974
rect 25975 10940 26000 10974
rect 25822 10867 25856 10901
rect 25894 10867 25928 10901
rect 25966 10867 25975 10901
rect 25975 10867 26000 10901
rect 25822 10794 25856 10828
rect 25894 10794 25928 10828
rect 25966 10794 25975 10828
rect 25975 10794 26000 10828
rect 25822 10721 25856 10755
rect 25894 10721 25928 10755
rect 25966 10721 25975 10755
rect 25975 10721 26000 10755
rect 25822 10648 25856 10682
rect 25894 10648 25928 10682
rect 25966 10648 25975 10682
rect 25975 10648 26000 10682
rect 1301 10550 1335 10584
rect 1382 10550 1416 10584
rect 1462 10550 1496 10584
rect 1542 10550 1576 10584
rect 1622 10550 1656 10584
rect 1702 10550 1736 10584
rect 1782 10550 1816 10584
rect 1862 10550 1877 10584
rect 1877 10550 1896 10584
rect 1942 10550 1972 10584
rect 1972 10550 1976 10584
rect 25822 10575 25856 10609
rect 25894 10575 25928 10609
rect 25966 10575 25975 10609
rect 25975 10575 26000 10609
rect 25822 10502 25856 10536
rect 25894 10502 25928 10536
rect 25966 10502 25975 10536
rect 25975 10502 26000 10536
rect 1687 10483 1721 10499
rect 1687 10465 1721 10483
rect 1687 10415 1721 10426
rect 1687 10392 1721 10415
rect 1687 10347 1721 10352
rect 1687 10318 1721 10347
rect 1843 10143 1877 10149
rect 1843 10115 1877 10143
rect 1843 10075 1877 10077
rect 1843 10043 1877 10075
rect 1999 10483 2033 10499
rect 1999 10465 2033 10483
rect 1999 10415 2033 10426
rect 1999 10392 2033 10415
rect 1999 10347 2033 10352
rect 1999 10318 2033 10347
rect 25822 10429 25856 10463
rect 25894 10429 25928 10463
rect 25966 10429 25975 10463
rect 25975 10429 26000 10463
rect 25822 10356 25856 10390
rect 25894 10356 25928 10390
rect 25966 10356 25975 10390
rect 25975 10356 26000 10390
rect 25822 10283 25856 10317
rect 25894 10283 25928 10317
rect 25966 10283 25975 10317
rect 25975 10283 26000 10317
rect 25822 10210 25856 10244
rect 25894 10210 25928 10244
rect 25966 10210 25975 10244
rect 25975 10210 26000 10244
rect 25822 10137 25856 10171
rect 25894 10137 25928 10171
rect 25966 10137 25975 10171
rect 25975 10137 26000 10171
rect 25822 10064 25856 10098
rect 25894 10064 25928 10098
rect 25966 10064 25975 10098
rect 25975 10064 26000 10098
rect 25822 9991 25856 10025
rect 25894 9991 25928 10025
rect 25966 9991 25975 10025
rect 25975 9991 26000 10025
rect 25822 9918 25856 9952
rect 25894 9918 25928 9952
rect 25966 9918 25975 9952
rect 25975 9918 26000 9952
rect 25822 9845 25856 9879
rect 25894 9845 25928 9879
rect 25966 9845 25975 9879
rect 25975 9845 26000 9879
rect 1301 9754 1305 9788
rect 1305 9754 1335 9788
rect 1400 9754 1434 9788
rect 1499 9754 1529 9788
rect 1529 9754 1533 9788
rect 25822 9772 25856 9806
rect 25894 9772 25928 9806
rect 25966 9772 25975 9806
rect 25975 9772 26000 9806
rect 903 9638 1005 9710
rect 1043 9637 1073 9671
rect 1073 9637 1077 9671
rect 899 9565 903 9599
rect 903 9565 933 9599
rect 971 9565 1005 9599
rect 1043 9564 1073 9598
rect 1073 9564 1077 9598
rect 899 9492 903 9526
rect 903 9492 933 9526
rect 971 9492 1005 9526
rect 1043 9491 1073 9525
rect 1073 9491 1077 9525
rect 899 9419 903 9453
rect 903 9419 933 9453
rect 971 9419 1005 9453
rect 1043 9418 1073 9452
rect 1073 9418 1077 9452
rect 899 9346 903 9380
rect 903 9346 933 9380
rect 971 9346 1005 9380
rect 1043 9345 1073 9379
rect 1073 9345 1077 9379
rect 899 9273 903 9307
rect 903 9273 933 9307
rect 971 9273 1005 9307
rect 1043 9272 1073 9306
rect 1073 9272 1077 9306
rect 899 9200 903 9234
rect 903 9200 933 9234
rect 971 9200 1005 9234
rect 1043 9199 1073 9233
rect 1073 9199 1077 9233
rect 899 9127 903 9161
rect 903 9127 933 9161
rect 971 9127 1005 9161
rect 1244 9687 1278 9691
rect 1244 9657 1278 9687
rect 1244 9585 1278 9618
rect 1244 9584 1278 9585
rect 1244 9517 1278 9544
rect 1244 9510 1278 9517
rect 1400 9449 1434 9454
rect 1400 9420 1434 9449
rect 1400 9381 1434 9382
rect 1400 9348 1434 9381
rect 1556 9687 1590 9691
rect 1556 9657 1590 9687
rect 1556 9585 1590 9618
rect 1556 9584 1590 9585
rect 1556 9517 1590 9544
rect 1556 9510 1590 9517
rect 25822 9699 25856 9733
rect 25894 9699 25928 9733
rect 25966 9699 25975 9733
rect 25975 9699 26000 9733
rect 25822 9626 25856 9660
rect 25894 9626 25928 9660
rect 25966 9626 25975 9660
rect 25975 9626 26000 9660
rect 25822 9553 25856 9587
rect 25894 9553 25928 9587
rect 25966 9553 25975 9587
rect 25975 9553 26000 9587
rect 25822 9480 25856 9514
rect 25894 9480 25928 9514
rect 25966 9480 25975 9514
rect 25975 9480 26000 9514
rect 25822 9407 25856 9441
rect 25894 9407 25928 9441
rect 25966 9407 25975 9441
rect 25975 9407 26000 9441
rect 25822 9334 25856 9368
rect 25894 9334 25928 9368
rect 25966 9334 25975 9368
rect 25975 9334 26000 9368
rect 25822 9261 25856 9295
rect 25894 9261 25928 9295
rect 25966 9261 25975 9295
rect 25975 9261 26000 9295
rect 25822 9188 25856 9222
rect 25894 9188 25928 9222
rect 25966 9188 25975 9222
rect 25975 9188 26000 9222
rect 1043 9126 1073 9160
rect 1073 9126 1077 9160
rect 899 9054 903 9088
rect 903 9054 933 9088
rect 971 9054 1005 9088
rect 1043 9053 1073 9087
rect 1073 9053 1077 9087
rect 899 8981 903 9015
rect 903 8981 933 9015
rect 971 8981 1005 9015
rect 1043 8980 1073 9014
rect 1073 8980 1077 9014
rect 899 8908 903 8942
rect 903 8908 933 8942
rect 971 8908 1005 8942
rect 1043 8907 1073 8941
rect 1073 8907 1077 8941
rect 899 8835 903 8869
rect 903 8835 933 8869
rect 971 8835 1005 8869
rect 1043 8834 1073 8868
rect 1073 8834 1077 8868
rect 899 8762 903 8796
rect 903 8762 933 8796
rect 971 8762 1005 8796
rect 1043 8761 1073 8795
rect 1073 8761 1077 8795
rect 899 8689 903 8723
rect 903 8689 933 8723
rect 971 8689 1005 8723
rect 1043 8688 1073 8722
rect 1073 8688 1077 8722
rect 899 8616 903 8650
rect 903 8616 933 8650
rect 971 8616 1005 8650
rect 1043 8615 1073 8649
rect 1073 8615 1077 8649
rect 899 8543 903 8577
rect 903 8543 933 8577
rect 971 8543 1005 8577
rect 1043 8542 1073 8576
rect 1073 8542 1077 8576
rect 899 8470 903 8504
rect 903 8470 933 8504
rect 971 8470 1005 8504
rect 1043 8469 1073 8503
rect 1073 8469 1077 8503
rect 899 8397 903 8431
rect 903 8397 933 8431
rect 971 8397 1005 8431
rect 1043 8396 1073 8430
rect 1073 8396 1077 8430
rect 899 8324 903 8358
rect 903 8324 933 8358
rect 971 8324 1005 8358
rect 1043 8323 1073 8357
rect 1073 8323 1077 8357
rect 899 8251 903 8285
rect 903 8251 933 8285
rect 971 8251 1005 8285
rect 1043 8250 1073 8284
rect 1073 8250 1077 8284
rect 899 8178 903 8212
rect 903 8178 933 8212
rect 971 8178 1005 8212
rect 1043 8177 1073 8211
rect 1073 8177 1077 8211
rect 899 8105 903 8139
rect 903 8105 933 8139
rect 971 8105 1005 8139
rect 25822 9115 25856 9149
rect 25894 9115 25928 9149
rect 25966 9115 25975 9149
rect 25975 9115 26000 9149
rect 25822 9042 25856 9076
rect 25894 9042 25928 9076
rect 25966 9042 25975 9076
rect 25975 9042 26000 9076
rect 25822 8969 25856 9003
rect 25894 8969 25928 9003
rect 25966 8969 25975 9003
rect 25975 8969 26000 9003
rect 25822 8896 25856 8930
rect 25894 8896 25928 8930
rect 25966 8896 25975 8930
rect 25975 8896 26000 8930
rect 25822 8823 25856 8857
rect 25894 8823 25928 8857
rect 25966 8823 25975 8857
rect 25975 8823 26000 8857
rect 25822 8750 25856 8784
rect 25894 8750 25928 8784
rect 25966 8750 25975 8784
rect 25975 8750 26000 8784
rect 25822 8677 25856 8711
rect 25894 8677 25928 8711
rect 25966 8677 25975 8711
rect 25975 8677 26000 8711
rect 25822 8604 25856 8638
rect 25894 8604 25928 8638
rect 25966 8604 25975 8638
rect 25975 8604 26000 8638
rect 25822 8531 25856 8565
rect 25894 8531 25928 8565
rect 25966 8531 25975 8565
rect 25975 8531 26000 8565
rect 25822 8458 25856 8492
rect 25894 8458 25928 8492
rect 25966 8458 25975 8492
rect 25975 8458 26000 8492
rect 25822 8385 25856 8419
rect 25894 8385 25928 8419
rect 25966 8385 25975 8419
rect 25975 8385 26000 8419
rect 25822 8312 25856 8346
rect 25894 8312 25928 8346
rect 25966 8312 25975 8346
rect 25975 8312 26000 8346
rect 25822 8239 25856 8273
rect 25894 8239 25928 8273
rect 25966 8239 25975 8273
rect 25975 8239 26000 8273
rect 1043 8104 1073 8138
rect 1073 8104 1077 8138
rect 25822 8166 25856 8200
rect 25894 8166 25928 8200
rect 25966 8166 25975 8200
rect 25975 8166 26000 8200
rect 899 8032 903 8066
rect 903 8032 933 8066
rect 971 8032 1005 8066
rect 1043 8031 1073 8065
rect 1073 8031 1077 8065
rect 899 7959 903 7993
rect 903 7959 933 7993
rect 971 7959 1005 7993
rect 1043 7958 1073 7992
rect 1073 7958 1077 7992
rect 899 7886 903 7920
rect 903 7886 933 7920
rect 971 7886 1005 7920
rect 1043 7885 1073 7919
rect 1073 7885 1077 7919
rect 899 7813 903 7847
rect 903 7813 933 7847
rect 971 7813 1005 7847
rect 1043 7812 1073 7846
rect 1073 7812 1077 7846
rect 899 7740 903 7774
rect 903 7740 933 7774
rect 971 7740 1005 7774
rect 1043 7739 1073 7773
rect 1073 7739 1077 7773
rect 899 7667 903 7701
rect 903 7667 933 7701
rect 971 7667 1005 7701
rect 1043 7666 1073 7700
rect 1073 7666 1077 7700
rect 899 7594 903 7628
rect 903 7594 933 7628
rect 971 7594 1005 7628
rect 1043 7593 1073 7627
rect 1073 7593 1077 7627
rect 899 7521 903 7555
rect 903 7521 933 7555
rect 971 7521 1005 7555
rect 1043 7520 1073 7554
rect 1073 7520 1077 7554
rect 899 7448 903 7482
rect 903 7448 933 7482
rect 971 7448 1005 7482
rect 1043 7447 1073 7481
rect 1073 7447 1077 7481
rect 899 7375 903 7409
rect 903 7375 933 7409
rect 971 7375 1005 7409
rect 1043 7374 1073 7408
rect 1073 7374 1077 7408
rect 899 7302 903 7336
rect 903 7302 933 7336
rect 971 7302 1005 7336
rect 1043 7301 1073 7335
rect 1073 7301 1077 7335
rect 899 7229 933 7263
rect 971 7229 1005 7263
rect 1043 7228 1077 7262
rect 899 7169 933 7190
rect 971 7169 1005 7190
rect 1043 7169 1077 7189
rect 899 7156 903 7169
rect 903 7156 933 7169
rect 971 7156 1005 7169
rect 1043 7155 1073 7169
rect 1073 7155 1077 7169
rect 899 7083 903 7117
rect 903 7083 933 7117
rect 971 7083 1005 7117
rect 1043 7082 1073 7116
rect 1073 7082 1077 7116
rect 899 7010 903 7044
rect 903 7010 933 7044
rect 971 7010 1005 7044
rect 1043 7009 1073 7043
rect 1073 7009 1077 7043
rect 899 6937 903 6971
rect 903 6937 933 6971
rect 971 6937 1005 6971
rect 1043 6936 1073 6970
rect 1073 6936 1077 6970
rect 899 6864 903 6898
rect 903 6864 933 6898
rect 971 6864 1005 6898
rect 1043 6863 1073 6897
rect 1073 6863 1077 6897
rect 25822 8093 25856 8127
rect 25894 8093 25928 8127
rect 25966 8093 25975 8127
rect 25975 8093 26000 8127
rect 25822 8020 25856 8054
rect 25894 8020 25928 8054
rect 25966 8020 25975 8054
rect 25975 8020 26000 8054
rect 25822 7947 25856 7981
rect 25894 7947 25928 7981
rect 25966 7947 25975 7981
rect 25975 7947 26000 7981
rect 25822 7874 25856 7908
rect 25894 7874 25928 7908
rect 25966 7874 25975 7908
rect 25975 7874 26000 7908
rect 25822 7801 25856 7835
rect 25894 7801 25928 7835
rect 25966 7801 25975 7835
rect 25975 7801 26000 7835
rect 25822 7728 25856 7762
rect 25894 7728 25928 7762
rect 25966 7728 25975 7762
rect 25975 7728 26000 7762
rect 25822 7655 25856 7689
rect 25894 7655 25928 7689
rect 25966 7655 25975 7689
rect 25975 7655 26000 7689
rect 899 6795 903 6825
rect 903 6795 933 6825
rect 971 6795 1005 6825
rect 1043 6820 25053 6824
rect 25092 6820 25126 6824
rect 25165 6820 25199 6824
rect 25238 6820 25272 6824
rect 25311 6820 25345 6824
rect 25384 6820 25418 6824
rect 25457 6820 25491 6824
rect 25530 6820 25564 6824
rect 25603 6820 25637 6824
rect 25676 6820 25710 6824
rect 25749 6820 25783 6824
rect 899 6791 933 6795
rect 971 6791 1005 6795
rect 1043 6752 25053 6820
rect 25092 6790 25126 6820
rect 25165 6790 25199 6820
rect 25238 6790 25272 6820
rect 25311 6790 25345 6820
rect 25384 6790 25418 6820
rect 25457 6790 25491 6820
rect 25530 6790 25564 6820
rect 25603 6790 25637 6820
rect 25676 6790 25710 6820
rect 25749 6790 25757 6820
rect 25757 6790 25783 6820
rect 25822 6790 25975 7616
rect 899 6727 903 6752
rect 903 6727 933 6752
rect 899 6718 933 6727
rect 971 6650 25125 6752
rect 25164 6718 25198 6752
rect 25237 6718 25271 6752
rect 25310 6718 25344 6752
rect 25383 6718 25417 6752
rect 25456 6718 25490 6752
rect 25529 6718 25563 6752
rect 25602 6718 25636 6752
rect 25675 6718 25709 6752
rect 25748 6718 25782 6752
rect 25821 6718 25825 6752
rect 25825 6718 25855 6752
rect 25894 6718 25975 6790
rect 25975 6718 26000 7616
rect 25164 6650 25198 6680
rect 25237 6650 25271 6680
rect 25310 6650 25344 6680
rect 25383 6650 25417 6680
rect 25456 6650 25490 6680
rect 25529 6650 25563 6680
rect 25602 6650 25636 6680
rect 25675 6650 25709 6680
rect 25748 6650 25782 6680
rect 25821 6650 25825 6680
rect 25825 6650 25855 6680
rect 971 6646 25125 6650
rect 25164 6646 25198 6650
rect 25237 6646 25271 6650
rect 25310 6646 25344 6650
rect 25383 6646 25417 6650
rect 25456 6646 25490 6650
rect 25529 6646 25563 6650
rect 25602 6646 25636 6650
rect 25675 6646 25709 6650
rect 25748 6646 25782 6650
rect 25821 6646 25855 6650
rect 25894 6646 25928 6680
rect 26220 12826 26224 12860
rect 26224 12826 26254 12860
rect 26292 12824 26326 12858
rect 26364 12824 26394 12858
rect 26394 12824 26398 12858
rect 26220 12752 26224 12786
rect 26224 12752 26254 12786
rect 26292 12750 26326 12784
rect 26364 12750 26394 12784
rect 26394 12750 26398 12784
rect 26220 12678 26224 12712
rect 26224 12678 26254 12712
rect 26292 12677 26326 12711
rect 26364 12677 26394 12711
rect 26394 12677 26398 12711
rect 26220 12604 26224 12638
rect 26224 12604 26254 12638
rect 26292 12604 26326 12638
rect 26364 12604 26394 12638
rect 26394 12604 26398 12638
rect 26220 12494 26224 12528
rect 26224 12494 26254 12528
rect 26292 12494 26326 12528
rect 26364 12494 26394 12528
rect 26394 12494 26398 12528
rect 26220 12421 26224 12455
rect 26224 12421 26254 12455
rect 26292 12421 26326 12455
rect 26364 12421 26394 12455
rect 26394 12421 26398 12455
rect 26220 12348 26224 12382
rect 26224 12348 26254 12382
rect 26292 12348 26326 12382
rect 26364 12348 26394 12382
rect 26394 12348 26398 12382
rect 26220 12275 26224 12309
rect 26224 12275 26254 12309
rect 26292 12275 26326 12309
rect 26364 12275 26394 12309
rect 26394 12275 26398 12309
rect 26220 12202 26224 12236
rect 26224 12202 26254 12236
rect 26292 12202 26326 12236
rect 26364 12202 26394 12236
rect 26394 12202 26398 12236
rect 657 6596 687 6630
rect 687 6596 691 6630
rect 513 6524 517 6558
rect 517 6524 547 6558
rect 585 6524 619 6558
rect 657 6523 687 6557
rect 687 6523 691 6557
rect 513 6451 517 6485
rect 517 6451 547 6485
rect 585 6451 619 6485
rect 657 6450 687 6484
rect 687 6450 691 6484
rect 513 6378 517 6412
rect 517 6378 547 6412
rect 585 6378 619 6412
rect 657 6377 687 6411
rect 687 6377 691 6411
rect 513 6305 517 6339
rect 517 6305 547 6339
rect 585 6305 619 6339
rect 657 6304 687 6338
rect 687 6304 691 6338
rect 513 6232 517 6266
rect 517 6232 547 6266
rect 585 6232 619 6266
rect 657 6231 687 6265
rect 687 6231 691 6265
rect 513 6159 517 6193
rect 517 6159 547 6193
rect 585 6159 619 6193
rect 657 6158 687 6192
rect 687 6158 691 6192
rect 513 6086 517 6120
rect 517 6086 547 6120
rect 585 6086 619 6120
rect 657 6085 687 6119
rect 687 6085 691 6119
rect 513 6013 517 6047
rect 517 6013 547 6047
rect 585 6013 619 6047
rect 657 6012 687 6046
rect 687 6012 691 6046
rect 513 5940 517 5974
rect 517 5940 547 5974
rect 585 5940 619 5974
rect 657 5939 687 5973
rect 687 5939 691 5973
rect 513 5867 517 5901
rect 517 5867 547 5901
rect 585 5867 619 5901
rect 657 5866 687 5900
rect 687 5866 691 5900
rect 26220 7680 26224 12163
rect 26224 7680 26394 12163
rect 26220 7645 26292 7680
rect 26220 7611 26224 7645
rect 26224 7611 26258 7645
rect 26258 7612 26292 7645
rect 26292 7612 26394 7680
rect 26394 7612 26398 12163
rect 26258 7611 26398 7612
rect 26220 7577 26398 7611
rect 26220 7576 26292 7577
rect 26220 7542 26224 7576
rect 26224 7542 26258 7576
rect 26258 7543 26292 7576
rect 26292 7543 26326 7577
rect 26326 7543 26360 7577
rect 26360 7543 26394 7577
rect 26394 7543 26398 7577
rect 26258 7542 26398 7543
rect 26220 7508 26398 7542
rect 26220 7507 26292 7508
rect 26220 7473 26224 7507
rect 26224 7473 26258 7507
rect 26258 7474 26292 7507
rect 26292 7474 26326 7508
rect 26326 7474 26360 7508
rect 26360 7474 26394 7508
rect 26394 7474 26398 7508
rect 26258 7473 26398 7474
rect 26220 7439 26398 7473
rect 26220 7438 26292 7439
rect 26220 7404 26224 7438
rect 26224 7404 26258 7438
rect 26258 7405 26292 7438
rect 26292 7405 26326 7439
rect 26326 7405 26360 7439
rect 26360 7405 26394 7439
rect 26394 7405 26398 7439
rect 26258 7404 26398 7405
rect 26220 7370 26398 7404
rect 26220 7369 26292 7370
rect 26220 7335 26224 7369
rect 26224 7335 26258 7369
rect 26258 7336 26292 7369
rect 26292 7336 26326 7370
rect 26326 7336 26360 7370
rect 26360 7336 26394 7370
rect 26394 7336 26398 7370
rect 26258 7335 26398 7336
rect 26220 7301 26398 7335
rect 26220 7300 26292 7301
rect 26220 7266 26224 7300
rect 26224 7266 26258 7300
rect 26258 7267 26292 7300
rect 26292 7267 26326 7301
rect 26326 7267 26360 7301
rect 26360 7267 26394 7301
rect 26394 7267 26398 7301
rect 26258 7266 26398 7267
rect 26220 7232 26398 7266
rect 26220 7231 26292 7232
rect 26220 7197 26224 7231
rect 26224 7197 26258 7231
rect 26258 7198 26292 7231
rect 26292 7198 26326 7232
rect 26326 7198 26360 7232
rect 26360 7198 26394 7232
rect 26394 7198 26398 7232
rect 26258 7197 26398 7198
rect 26220 7163 26398 7197
rect 26220 7162 26292 7163
rect 26220 7128 26224 7162
rect 26224 7128 26258 7162
rect 26258 7129 26292 7162
rect 26292 7129 26326 7163
rect 26326 7129 26360 7163
rect 26360 7129 26394 7163
rect 26394 7129 26398 7163
rect 26258 7128 26398 7129
rect 26220 7094 26398 7128
rect 26220 7093 26292 7094
rect 26220 7059 26224 7093
rect 26224 7059 26258 7093
rect 26258 7060 26292 7093
rect 26292 7060 26326 7094
rect 26326 7060 26360 7094
rect 26360 7060 26394 7094
rect 26394 7060 26398 7094
rect 26258 7059 26398 7060
rect 26220 7025 26398 7059
rect 26220 7024 26292 7025
rect 26220 6990 26224 7024
rect 26224 6990 26258 7024
rect 26258 6991 26292 7024
rect 26292 6991 26326 7025
rect 26326 6991 26360 7025
rect 26360 6991 26394 7025
rect 26394 6991 26398 7025
rect 26258 6990 26398 6991
rect 26220 6956 26398 6990
rect 26220 6955 26292 6956
rect 26220 6921 26224 6955
rect 26224 6921 26258 6955
rect 26258 6922 26292 6955
rect 26292 6922 26326 6956
rect 26326 6922 26360 6956
rect 26360 6922 26394 6956
rect 26394 6922 26398 6956
rect 26258 6921 26398 6922
rect 26220 6887 26398 6921
rect 26220 6886 26292 6887
rect 26220 6852 26224 6886
rect 26224 6852 26258 6886
rect 26258 6853 26292 6886
rect 26292 6853 26326 6887
rect 26326 6853 26360 6887
rect 26360 6853 26394 6887
rect 26394 6853 26398 6887
rect 26258 6852 26398 6853
rect 26220 6818 26398 6852
rect 26220 6817 26292 6818
rect 26220 6783 26224 6817
rect 26224 6783 26258 6817
rect 26258 6784 26292 6817
rect 26292 6784 26326 6818
rect 26326 6784 26360 6818
rect 26360 6784 26394 6818
rect 26394 6784 26398 6818
rect 26258 6783 26398 6784
rect 26220 6749 26398 6783
rect 26220 6748 26292 6749
rect 26220 6714 26224 6748
rect 26224 6714 26258 6748
rect 26258 6715 26292 6748
rect 26292 6715 26326 6749
rect 26326 6715 26360 6749
rect 26360 6715 26394 6749
rect 26394 6715 26398 6749
rect 26258 6714 26398 6715
rect 26220 6680 26398 6714
rect 26220 6679 26292 6680
rect 26220 6645 26224 6679
rect 26224 6645 26258 6679
rect 26258 6646 26292 6679
rect 26292 6646 26326 6680
rect 26326 6646 26360 6680
rect 26360 6646 26394 6680
rect 26394 6646 26398 6680
rect 26258 6645 26398 6646
rect 26220 6611 26398 6645
rect 26220 6610 26292 6611
rect 26220 6576 26224 6610
rect 26224 6576 26258 6610
rect 26258 6577 26292 6610
rect 26292 6577 26326 6611
rect 26326 6577 26360 6611
rect 26360 6577 26394 6611
rect 26394 6577 26398 6611
rect 26258 6576 26398 6577
rect 26220 6542 26398 6576
rect 26220 6541 26292 6542
rect 26220 6507 26224 6541
rect 26224 6507 26258 6541
rect 26258 6508 26292 6541
rect 26292 6508 26326 6542
rect 26326 6508 26360 6542
rect 26360 6508 26394 6542
rect 26394 6508 26398 6542
rect 26258 6507 26398 6508
rect 26220 6473 26398 6507
rect 26220 6472 26292 6473
rect 26220 6438 26224 6472
rect 26224 6438 26258 6472
rect 26258 6439 26292 6472
rect 26292 6439 26326 6473
rect 26326 6439 26360 6473
rect 26360 6439 26394 6473
rect 26394 6439 26398 6473
rect 26258 6438 26398 6439
rect 26220 6404 26398 6438
rect 26220 6403 26292 6404
rect 26220 6369 26224 6403
rect 26224 6369 26258 6403
rect 26258 6370 26292 6403
rect 26292 6370 26326 6404
rect 26326 6370 26360 6404
rect 26360 6370 26394 6404
rect 26394 6370 26398 6404
rect 26258 6369 26398 6370
rect 26220 6335 26398 6369
rect 26220 6334 26292 6335
rect 26220 6300 26224 6334
rect 26224 6300 26258 6334
rect 26258 6301 26292 6334
rect 26292 6301 26326 6335
rect 26326 6301 26360 6335
rect 26360 6301 26394 6335
rect 26394 6301 26398 6335
rect 26258 6300 26398 6301
rect 26220 6266 26398 6300
rect 26220 6265 26292 6266
rect 26220 6231 26224 6265
rect 26224 6231 26258 6265
rect 26258 6232 26292 6265
rect 26292 6232 26326 6266
rect 26326 6232 26360 6266
rect 26360 6232 26394 6266
rect 26394 6232 26398 6266
rect 26258 6231 26398 6232
rect 26220 6197 26398 6231
rect 26220 6196 26292 6197
rect 26220 6162 26224 6196
rect 26224 6162 26258 6196
rect 26258 6163 26292 6196
rect 26292 6163 26326 6197
rect 26326 6163 26360 6197
rect 26360 6163 26394 6197
rect 26394 6163 26398 6197
rect 26258 6162 26398 6163
rect 26220 6128 26398 6162
rect 26220 6127 26292 6128
rect 26220 6093 26224 6127
rect 26224 6093 26258 6127
rect 26258 6094 26292 6127
rect 26292 6094 26326 6128
rect 26326 6094 26360 6128
rect 26360 6094 26394 6128
rect 26394 6094 26398 6128
rect 26258 6093 26398 6094
rect 26220 6059 26398 6093
rect 26220 6058 26292 6059
rect 26220 6024 26224 6058
rect 26224 6024 26258 6058
rect 26258 6025 26292 6058
rect 26292 6025 26326 6059
rect 26326 6025 26360 6059
rect 26360 6025 26394 6059
rect 26394 6025 26398 6059
rect 26258 6024 26398 6025
rect 26220 5990 26398 6024
rect 26220 5989 26292 5990
rect 26220 5955 26224 5989
rect 26224 5955 26258 5989
rect 26258 5956 26292 5989
rect 26292 5956 26326 5990
rect 26326 5956 26360 5990
rect 26360 5956 26394 5990
rect 26394 5956 26398 5990
rect 26258 5955 26398 5956
rect 26220 5921 26398 5955
rect 26220 5920 26292 5921
rect 26220 5886 26224 5920
rect 26224 5886 26258 5920
rect 26258 5887 26292 5920
rect 26292 5887 26326 5921
rect 26326 5887 26360 5921
rect 26360 5887 26394 5921
rect 26394 5887 26398 5921
rect 26258 5886 26398 5887
rect 26220 5852 26398 5886
rect 26220 5851 26292 5852
rect 513 5794 517 5828
rect 517 5794 547 5828
rect 585 5794 619 5828
rect 657 5817 687 5827
rect 687 5817 722 5827
rect 722 5817 756 5827
rect 756 5817 791 5827
rect 791 5817 825 5827
rect 825 5817 860 5827
rect 657 5783 860 5817
rect 860 5783 26035 5827
rect 26074 5793 26108 5827
rect 26147 5793 26181 5827
rect 26220 5793 26258 5851
rect 26258 5818 26292 5851
rect 26292 5818 26326 5852
rect 26326 5818 26360 5852
rect 26360 5818 26394 5852
rect 26394 5818 26398 5852
rect 26258 5793 26398 5818
rect 26292 5783 26398 5793
rect 657 5755 688 5783
rect 513 5749 517 5755
rect 517 5749 547 5755
rect 585 5749 619 5755
rect 619 5749 654 5755
rect 654 5749 688 5755
rect 688 5749 723 5783
rect 723 5749 757 5783
rect 757 5749 792 5783
rect 792 5755 26035 5783
rect 513 5721 547 5749
rect 585 5715 792 5749
rect 585 5681 619 5715
rect 619 5681 654 5715
rect 654 5681 688 5715
rect 688 5681 723 5715
rect 723 5681 757 5715
rect 757 5681 792 5715
rect 792 5681 26107 5755
rect 26146 5721 26180 5755
rect 26219 5721 26253 5755
rect 26292 5721 26326 5783
rect 26326 5749 26360 5783
rect 26360 5749 26394 5783
rect 26394 5749 26398 5783
rect 26326 5721 26398 5749
rect 26146 5681 26180 5683
rect 26219 5681 26253 5683
rect 26292 5681 26326 5683
rect 585 5649 26107 5681
rect 26146 5649 26180 5681
rect 26219 5649 26253 5681
rect 26292 5649 26326 5681
rect -619 3032 -585 3066
rect -533 3032 -499 3066
rect -447 3032 -413 3066
rect -362 3032 -328 3066
rect -277 3032 -243 3066
rect -619 2954 -585 2988
rect -533 2954 -499 2988
rect -447 2954 -413 2988
rect -362 2954 -328 2988
rect -277 2954 -243 2988
rect -139 3032 -105 3066
rect -53 3032 -19 3066
rect 33 3032 67 3066
rect 118 3032 152 3066
rect 203 3032 237 3066
rect -139 2954 -105 2988
rect -53 2954 -19 2988
rect 33 2954 67 2988
rect 118 2954 152 2988
rect 203 2954 237 2988
rect 346 3032 380 3066
rect 432 3032 466 3066
rect 518 3032 552 3066
rect 603 3032 637 3066
rect 688 3032 722 3066
rect 346 2954 380 2988
rect 432 2954 466 2988
rect 518 2954 552 2988
rect 603 2954 637 2988
rect 688 2954 722 2988
rect -1123 2892 -1089 2926
rect -1035 2892 -1001 2926
rect -948 2892 -914 2926
rect -861 2892 -827 2926
rect -774 2892 -740 2926
rect 24517 3017 24551 3033
rect 24517 2999 24551 3017
rect 24517 2915 24551 2933
rect 24517 2899 24551 2915
rect -1123 2806 -1089 2840
rect -1035 2806 -1001 2840
rect -948 2806 -914 2840
rect -861 2806 -827 2840
rect -774 2806 -740 2840
rect 24517 2699 24551 2715
rect 24517 2681 24551 2699
rect 24517 2631 24551 2643
rect 24517 2609 24551 2631
rect -1132 1260 -1098 1294
rect -1058 1260 -1024 1294
rect -984 1260 -950 1294
rect -910 1260 -876 1294
rect -836 1260 -802 1294
rect -762 1260 -728 1294
rect -688 1260 -654 1294
rect -614 1260 -580 1294
rect -540 1260 -506 1294
rect -466 1260 -432 1294
rect -392 1260 -358 1294
rect -319 1260 -285 1294
rect -246 1260 -212 1294
rect -173 1260 -139 1294
rect -100 1260 -66 1294
rect -27 1260 7 1294
rect 46 1260 80 1294
rect 119 1260 153 1294
rect 192 1260 226 1294
rect 265 1260 299 1294
rect 338 1260 372 1294
rect 411 1260 445 1294
rect 484 1260 518 1294
rect 557 1260 591 1294
rect 630 1260 664 1294
rect 703 1260 737 1294
rect -1132 1186 -1098 1220
rect -1058 1186 -1024 1220
rect -984 1186 -950 1220
rect -910 1186 -876 1220
rect -836 1186 -802 1220
rect -762 1186 -728 1220
rect -688 1186 -654 1220
rect -614 1186 -580 1220
rect -540 1186 -506 1220
rect -466 1186 -432 1220
rect -392 1186 -358 1220
rect -319 1186 -285 1220
rect -246 1186 -212 1220
rect -173 1186 -139 1220
rect -100 1186 -66 1220
rect -27 1186 7 1220
rect 46 1186 80 1220
rect 119 1186 153 1220
rect 192 1186 226 1220
rect 265 1186 299 1220
rect 338 1186 372 1220
rect 411 1186 445 1220
rect 484 1186 518 1220
rect 557 1186 591 1220
rect 630 1186 664 1220
rect 703 1186 737 1220
rect -1132 1112 -1098 1146
rect -1058 1112 -1024 1146
rect -984 1112 -950 1146
rect -910 1112 -876 1146
rect -836 1112 -802 1146
rect -762 1112 -728 1146
rect -688 1112 -654 1146
rect -614 1112 -580 1146
rect -540 1112 -506 1146
rect -466 1112 -432 1146
rect -392 1112 -358 1146
rect -319 1112 -285 1146
rect -246 1112 -212 1146
rect -173 1112 -139 1146
rect -100 1112 -66 1146
rect -27 1112 7 1146
rect 46 1112 80 1146
rect 119 1112 153 1146
rect 192 1112 226 1146
rect 265 1112 299 1146
rect 338 1112 372 1146
rect 411 1112 445 1146
rect 484 1112 518 1146
rect 557 1112 591 1146
rect 630 1112 664 1146
rect 703 1112 737 1146
rect -1132 1038 -1098 1072
rect -1058 1038 -1024 1072
rect -984 1038 -950 1072
rect -910 1038 -876 1072
rect -836 1038 -802 1072
rect -762 1038 -728 1072
rect -688 1038 -654 1072
rect -614 1038 -580 1072
rect -540 1038 -506 1072
rect -466 1038 -432 1072
rect -392 1038 -358 1072
rect -319 1038 -285 1072
rect -246 1038 -212 1072
rect -173 1038 -139 1072
rect -100 1038 -66 1072
rect -27 1038 7 1072
rect 46 1038 80 1072
rect 119 1038 153 1072
rect 192 1038 226 1072
rect 265 1038 299 1072
rect 338 1038 372 1072
rect 411 1038 445 1072
rect 484 1038 518 1072
rect 557 1038 591 1072
rect 630 1038 664 1072
rect 703 1038 737 1072
rect -1132 964 -1098 998
rect -1058 964 -1024 998
rect -984 964 -950 998
rect -910 964 -876 998
rect -836 964 -802 998
rect -762 964 -728 998
rect -688 964 -654 998
rect -614 964 -580 998
rect -540 964 -506 998
rect -466 964 -432 998
rect -392 964 -358 998
rect -319 964 -285 998
rect -246 964 -212 998
rect -173 964 -139 998
rect -100 964 -66 998
rect -27 964 7 998
rect 46 964 80 998
rect 119 964 153 998
rect 192 964 226 998
rect 265 964 299 998
rect 338 964 372 998
rect 411 964 445 998
rect 484 964 518 998
rect 557 964 591 998
rect 630 964 664 998
rect 703 964 737 998
rect -1132 890 -1098 924
rect -1058 890 -1024 924
rect -984 890 -950 924
rect -910 890 -876 924
rect -836 890 -802 924
rect -762 890 -728 924
rect -688 890 -654 924
rect -614 890 -580 924
rect -540 890 -506 924
rect -466 890 -432 924
rect -392 890 -358 924
rect -319 890 -285 924
rect -246 890 -212 924
rect -173 890 -139 924
rect -100 890 -66 924
rect -27 890 7 924
rect 46 890 80 924
rect 119 890 153 924
rect 192 890 226 924
rect 265 890 299 924
rect 338 890 372 924
rect 411 890 445 924
rect 484 890 518 924
rect 557 890 591 924
rect 630 890 664 924
rect 703 890 737 924
rect -1132 816 -1098 850
rect -1058 816 -1024 850
rect -984 816 -950 850
rect -910 816 -876 850
rect -836 816 -802 850
rect -762 816 -728 850
rect -688 816 -654 850
rect -614 816 -580 850
rect -540 816 -506 850
rect -466 816 -432 850
rect -392 816 -358 850
rect -319 816 -285 850
rect -246 816 -212 850
rect -173 816 -139 850
rect -100 816 -66 850
rect -27 816 7 850
rect 46 816 80 850
rect 119 816 153 850
rect 192 816 226 850
rect 265 816 299 850
rect 338 816 372 850
rect 411 816 445 850
rect 484 816 518 850
rect 557 816 591 850
rect 630 816 664 850
rect 703 816 737 850
rect 23779 1159 23780 1193
rect 23780 1159 23813 1193
rect 23852 1159 23882 1193
rect 23882 1159 23886 1193
rect 23925 1159 23950 1193
rect 23950 1159 23959 1193
rect 23998 1159 24018 1193
rect 24018 1159 24032 1193
rect 24071 1159 24086 1193
rect 24086 1159 24105 1193
rect 24144 1159 24154 1193
rect 24154 1159 24178 1193
rect 24217 1159 24222 1193
rect 24222 1159 24251 1193
rect 24290 1159 24324 1193
rect 24363 1159 24392 1193
rect 24392 1159 24397 1193
rect 24436 1159 24460 1193
rect 24460 1159 24470 1193
rect 24509 1159 24528 1193
rect 24528 1159 24543 1193
rect 24582 1159 24596 1193
rect 24596 1159 24616 1193
rect 24655 1159 24664 1193
rect 24664 1159 24689 1193
rect 24728 1159 24732 1193
rect 24732 1159 24762 1193
rect 24801 1159 24834 1193
rect 24834 1159 24835 1193
rect 24874 1159 24902 1193
rect 24902 1159 24908 1193
rect 24947 1159 24970 1193
rect 24970 1159 24981 1193
rect 25020 1159 25038 1193
rect 25038 1159 25054 1193
rect 25093 1159 25106 1193
rect 25106 1159 25127 1193
rect 25166 1159 25174 1193
rect 25174 1159 25200 1193
rect 25239 1159 25242 1193
rect 25242 1159 25273 1193
rect 25312 1159 25344 1193
rect 25344 1159 25346 1193
rect 25385 1159 25412 1193
rect 25412 1159 25419 1193
rect 25458 1159 25480 1193
rect 25480 1159 25492 1193
rect 25531 1159 25548 1193
rect 25548 1159 25565 1193
rect 25604 1159 25616 1193
rect 25616 1159 25638 1193
rect 25676 1159 25684 1193
rect 25684 1159 25710 1193
rect 25748 1159 25752 1193
rect 25752 1159 25782 1193
rect 23707 1091 23741 1105
rect 23707 1071 23741 1091
rect 24426 1076 24460 1110
rect 24500 1076 24534 1110
rect 24574 1076 24608 1110
rect 24648 1076 24682 1110
rect 24130 1027 24164 1029
rect 24229 1027 24263 1029
rect 24328 1027 24362 1029
rect 25186 1076 25220 1110
rect 25260 1076 25294 1110
rect 25334 1076 25368 1110
rect 25408 1076 25442 1110
rect 24899 1027 24933 1029
rect 24992 1027 25026 1029
rect 25084 1027 25118 1029
rect 24130 995 24164 1027
rect 24229 995 24259 1027
rect 24259 995 24263 1027
rect 24328 995 24354 1027
rect 24354 995 24362 1027
rect 24899 995 24924 1027
rect 24924 995 24933 1027
rect 24992 995 25019 1027
rect 25019 995 25026 1027
rect 25084 995 25114 1027
rect 25114 995 25118 1027
rect 25820 1091 25854 1121
rect 25820 1087 25854 1091
rect 25820 1023 25854 1042
rect 25820 1008 25854 1023
rect 23707 955 23741 979
rect 23707 945 23741 955
rect 23707 887 23741 893
rect 23707 859 23741 887
rect 23953 919 23987 945
rect 23953 911 23987 919
rect 24056 933 24090 934
rect 24056 900 24069 933
rect 24069 900 24090 933
rect 24128 900 24162 934
rect 24347 900 24381 934
rect 23953 839 23987 873
rect 23707 785 23741 807
rect 23707 773 23741 785
rect 24419 900 24453 934
rect 25569 938 25603 972
rect 24630 900 24664 934
rect 24702 933 24736 934
rect 24702 900 24727 933
rect 24727 900 24736 933
rect 24215 802 24249 836
rect 24287 802 24321 836
rect 24477 802 24511 836
rect 24549 802 24583 836
rect 24829 873 24863 906
rect 24937 893 24971 927
rect 25009 907 25043 927
rect 25009 893 25019 907
rect 25019 893 25043 907
rect 24829 872 24863 873
rect 25107 859 25141 893
rect 25277 907 25311 927
rect 25277 893 25297 907
rect 25297 893 25311 907
rect 25349 893 25383 927
rect 25179 859 25213 893
rect 25453 873 25487 890
rect 24829 800 24863 834
rect 25453 856 25487 873
rect 25569 885 25603 900
rect 25569 866 25603 885
rect 25820 955 25854 963
rect 25820 929 25854 955
rect 25453 784 25487 818
rect 25820 853 25854 884
rect 25820 850 25854 853
rect 23707 687 23741 721
rect 25820 785 25854 805
rect 25820 771 25854 785
rect 25820 717 25854 727
rect 25820 693 25854 717
rect 23779 615 23809 649
rect 23809 615 23813 649
rect 23851 615 23877 649
rect 23877 615 23885 649
rect 23923 615 23945 649
rect 23945 615 23957 649
rect 23996 615 24013 649
rect 24013 615 24030 649
rect 24069 615 24081 649
rect 24081 615 24103 649
rect 24142 615 24149 649
rect 24149 615 24176 649
rect 24215 615 24217 649
rect 24217 615 24249 649
rect 24288 615 24319 649
rect 24319 615 24322 649
rect 24361 615 24387 649
rect 24387 615 24395 649
rect 24434 615 24455 649
rect 24455 615 24468 649
rect 24507 615 24523 649
rect 24523 615 24541 649
rect 24580 615 24591 649
rect 24591 615 24614 649
rect 24653 615 24659 649
rect 24659 615 24687 649
rect 24726 615 24727 649
rect 24727 615 24760 649
rect 24799 615 24829 649
rect 24829 615 24833 649
rect 24872 615 24897 649
rect 24897 615 24906 649
rect 24945 615 24965 649
rect 24965 615 24979 649
rect 25018 615 25033 649
rect 25033 615 25052 649
rect 25091 615 25101 649
rect 25101 615 25125 649
rect 25164 615 25169 649
rect 25169 615 25198 649
rect 25237 615 25271 649
rect 25310 615 25339 649
rect 25339 615 25344 649
rect 25383 615 25407 649
rect 25407 615 25417 649
rect 25456 615 25475 649
rect 25475 615 25490 649
rect 25529 615 25543 649
rect 25543 615 25563 649
rect 25602 615 25611 649
rect 25611 615 25636 649
rect 25675 615 25679 649
rect 25679 615 25709 649
rect 25748 615 25781 649
rect 25781 615 25782 649
<< metal1 >>
rect 1090 22667 1832 22673
rect 1090 22633 1174 22667
rect 1208 22633 1252 22667
rect 1286 22633 1330 22667
rect 1364 22633 1408 22667
rect 1442 22633 1486 22667
rect 1520 22633 1564 22667
rect 1598 22633 1642 22667
rect 1676 22633 1720 22667
rect 1754 22633 1832 22667
rect 1090 22595 1832 22633
rect 1090 22561 1096 22595
rect 1130 22561 1168 22595
rect 1202 22561 1252 22595
rect 1286 22561 1330 22595
rect 1364 22561 1408 22595
rect 1442 22561 1486 22595
rect 1520 22561 1564 22595
rect 1598 22561 1642 22595
rect 1676 22561 1720 22595
rect 1090 22555 1720 22561
rect 1090 22522 1208 22555
rect 1090 22488 1096 22522
rect 1130 22488 1168 22522
rect 1202 22488 1208 22522
rect 1090 22449 1208 22488
rect 1090 22415 1096 22449
rect 1130 22415 1168 22449
rect 1202 22415 1208 22449
rect 1090 22376 1208 22415
rect 1714 22489 1720 22555
rect 1826 22489 1832 22595
rect 1714 22450 1832 22489
rect 1714 22416 1720 22450
rect 1754 22416 1792 22450
rect 1826 22416 1832 22450
rect 1090 22342 1096 22376
rect 1130 22342 1168 22376
rect 1202 22342 1208 22376
rect 1090 22303 1208 22342
rect 1090 22269 1096 22303
rect 1130 22269 1168 22303
rect 1202 22269 1208 22303
rect 1357 22407 1409 22413
rect 1357 22343 1409 22355
rect 1357 22287 1366 22291
rect 1400 22287 1409 22291
rect 1357 22278 1409 22287
tri 1357 22275 1360 22278 ne
rect 1360 22275 1406 22278
tri 1406 22275 1409 22278 nw
rect 1513 22407 1565 22413
rect 1513 22343 1565 22355
rect 1513 22287 1522 22291
rect 1556 22287 1565 22291
rect 1513 22278 1565 22287
tri 1513 22275 1516 22278 ne
rect 1516 22275 1562 22278
tri 1562 22275 1565 22278 nw
rect 1714 22377 1832 22416
rect 1714 22343 1720 22377
rect 1754 22343 1792 22377
rect 1826 22343 1832 22377
rect 1714 22304 1832 22343
rect 1090 22230 1208 22269
rect 1714 22270 1720 22304
rect 1754 22270 1792 22304
rect 1826 22270 1832 22304
rect 1090 22196 1096 22230
rect 1130 22196 1168 22230
rect 1202 22196 1208 22230
rect 1090 22157 1208 22196
rect 1090 22123 1096 22157
rect 1130 22123 1168 22157
rect 1202 22123 1208 22157
rect 1090 22084 1208 22123
rect 1090 22050 1096 22084
rect 1130 22050 1168 22084
rect 1202 22050 1208 22084
rect 1090 22011 1208 22050
rect 1090 21977 1096 22011
rect 1130 21977 1168 22011
rect 1202 21977 1208 22011
rect 1090 21938 1208 21977
rect 1090 16432 1096 21938
rect 1202 16472 1208 21938
rect 1282 22255 1328 22267
rect 1282 22221 1288 22255
rect 1322 22221 1328 22255
rect 1282 22183 1328 22221
rect 1282 22149 1288 22183
rect 1322 22149 1328 22183
rect 1282 22111 1328 22149
rect 1282 22077 1288 22111
rect 1322 22077 1328 22111
rect 1282 22039 1328 22077
rect 1435 22255 1487 22267
rect 1435 22245 1444 22255
rect 1478 22245 1487 22255
rect 1435 22183 1487 22193
rect 1435 22181 1444 22183
rect 1478 22181 1487 22183
rect 1435 22117 1487 22129
rect 1435 22059 1487 22065
tri 1435 22056 1438 22059 ne
rect 1282 22005 1288 22039
rect 1322 22005 1328 22039
rect 1282 21967 1328 22005
rect 1282 21933 1288 21967
rect 1322 21933 1328 21967
tri 1279 21913 1282 21916 se
rect 1282 21913 1328 21933
rect 1438 22039 1484 22059
tri 1484 22056 1487 22059 nw
rect 1594 22255 1640 22267
rect 1594 22221 1600 22255
rect 1634 22221 1640 22255
rect 1594 22183 1640 22221
rect 1594 22149 1600 22183
rect 1634 22149 1640 22183
rect 1594 22111 1640 22149
rect 1594 22077 1600 22111
rect 1634 22077 1640 22111
rect 1438 22005 1444 22039
rect 1478 22005 1484 22039
rect 1438 21967 1484 22005
rect 1438 21933 1444 21967
rect 1478 21933 1484 21967
tri 1328 21913 1331 21916 sw
rect 1279 21907 1331 21913
rect 1279 21843 1331 21855
rect 1279 21789 1288 21791
rect 1322 21789 1331 21791
rect 1279 21779 1331 21789
rect 1279 21717 1288 21727
rect 1322 21717 1331 21727
rect 1438 21895 1484 21933
rect 1594 22039 1640 22077
rect 1594 22005 1600 22039
rect 1634 22005 1640 22039
rect 1594 21967 1640 22005
rect 1594 21933 1600 21967
rect 1634 21933 1640 21967
rect 1438 21861 1444 21895
rect 1478 21861 1484 21895
rect 1438 21823 1484 21861
rect 1438 21789 1444 21823
rect 1478 21789 1484 21823
rect 1438 21751 1484 21789
rect 1279 21705 1331 21717
rect 1360 21708 1406 21720
rect 1360 21674 1366 21708
rect 1400 21674 1406 21708
rect 1438 21717 1444 21751
rect 1478 21717 1484 21751
tri 1591 21913 1594 21916 se
rect 1594 21913 1640 21933
rect 1714 22231 1832 22270
rect 1714 22197 1720 22231
rect 1754 22197 1792 22231
rect 1826 22197 1832 22231
rect 1714 22158 1832 22197
rect 1714 22124 1720 22158
rect 1754 22124 1792 22158
rect 1826 22124 1832 22158
rect 1714 22085 1832 22124
rect 1714 22051 1720 22085
rect 1754 22051 1792 22085
rect 1826 22051 1832 22085
rect 1714 22012 1832 22051
rect 1714 21978 1720 22012
rect 1754 21978 1792 22012
rect 1826 21978 1832 22012
rect 1714 21939 1832 21978
tri 1640 21913 1643 21916 sw
rect 1591 21907 1643 21913
rect 1591 21843 1643 21855
rect 1591 21789 1600 21791
rect 1634 21789 1643 21791
rect 1591 21779 1643 21789
rect 1438 21705 1484 21717
rect 1516 21708 1562 21720
rect 1360 21636 1406 21674
rect 1279 21593 1331 21605
rect 1279 21583 1288 21593
rect 1322 21583 1331 21593
rect 1360 21602 1366 21636
rect 1400 21602 1406 21636
rect 1516 21674 1522 21708
rect 1556 21674 1562 21708
rect 1591 21717 1600 21727
rect 1634 21717 1643 21727
rect 1591 21705 1643 21717
rect 1714 21905 1720 21939
rect 1754 21905 1792 21939
rect 1826 21905 1832 21939
rect 1714 21866 1832 21905
rect 1714 21832 1720 21866
rect 1754 21832 1792 21866
rect 1826 21832 1832 21866
rect 1714 21793 1832 21832
rect 1714 21759 1720 21793
rect 1754 21759 1792 21793
rect 1826 21759 1832 21793
rect 1714 21720 1832 21759
rect 1516 21636 1562 21674
rect 1360 21590 1406 21602
rect 1438 21593 1484 21605
rect 1279 21521 1331 21531
rect 1279 21519 1288 21521
rect 1322 21519 1331 21521
rect 1279 21455 1331 21467
rect 1279 21397 1331 21403
tri 1279 21394 1282 21397 ne
rect 1282 21377 1328 21397
tri 1328 21394 1331 21397 nw
rect 1438 21559 1444 21593
rect 1478 21559 1484 21593
rect 1516 21602 1522 21636
rect 1556 21602 1562 21636
rect 1714 21686 1720 21720
rect 1754 21686 1792 21720
rect 1826 21686 1832 21720
rect 1714 21647 1832 21686
rect 1714 21613 1720 21647
rect 1754 21613 1792 21647
rect 1826 21613 1832 21647
rect 1516 21590 1562 21602
rect 1591 21593 1643 21605
rect 1438 21521 1484 21559
rect 1438 21487 1444 21521
rect 1478 21487 1484 21521
rect 1438 21449 1484 21487
rect 1438 21415 1444 21449
rect 1478 21415 1484 21449
rect 1282 21343 1288 21377
rect 1322 21343 1328 21377
rect 1282 21305 1328 21343
rect 1282 21271 1288 21305
rect 1322 21271 1328 21305
rect 1282 21233 1328 21271
rect 1438 21377 1484 21415
rect 1591 21583 1600 21593
rect 1634 21583 1643 21593
rect 1591 21521 1643 21531
rect 1591 21519 1600 21521
rect 1634 21519 1643 21521
rect 1591 21455 1643 21467
rect 1591 21397 1643 21403
tri 1591 21394 1594 21397 ne
rect 1438 21343 1444 21377
rect 1478 21343 1484 21377
rect 1438 21305 1484 21343
rect 1438 21271 1444 21305
rect 1478 21271 1484 21305
rect 1282 21199 1288 21233
rect 1322 21199 1328 21233
rect 1282 21161 1328 21199
rect 1282 21127 1288 21161
rect 1322 21127 1328 21161
rect 1282 21089 1328 21127
rect 1282 21055 1288 21089
rect 1322 21055 1328 21089
rect 1282 21043 1328 21055
tri 1435 21251 1438 21254 se
rect 1438 21251 1484 21271
rect 1594 21377 1640 21397
tri 1640 21394 1643 21397 nw
rect 1714 21574 1832 21613
rect 1714 21540 1720 21574
rect 1754 21540 1792 21574
rect 1826 21540 1832 21574
rect 1714 21501 1832 21540
rect 1714 21467 1720 21501
rect 1754 21467 1792 21501
rect 1826 21467 1832 21501
rect 1714 21428 1832 21467
rect 1714 21394 1720 21428
rect 1754 21394 1792 21428
rect 1826 21394 1832 21428
rect 1594 21343 1600 21377
rect 1634 21343 1640 21377
rect 1594 21305 1640 21343
rect 1594 21271 1600 21305
rect 1634 21271 1640 21305
tri 1484 21251 1487 21254 sw
rect 1435 21245 1487 21251
rect 1435 21181 1487 21193
rect 1435 21127 1444 21129
rect 1478 21127 1487 21129
rect 1435 21117 1487 21127
rect 1435 21055 1444 21065
rect 1478 21055 1487 21065
rect 1435 21043 1487 21055
rect 1594 21233 1640 21271
rect 1594 21199 1600 21233
rect 1634 21199 1640 21233
rect 1594 21161 1640 21199
rect 1594 21127 1600 21161
rect 1634 21127 1640 21161
rect 1594 21089 1640 21127
rect 1594 21055 1600 21089
rect 1634 21055 1640 21089
rect 1714 21355 1832 21394
rect 1714 21321 1720 21355
rect 1754 21321 1792 21355
rect 1826 21321 1832 21355
rect 1714 21282 1832 21321
rect 1714 21248 1720 21282
rect 1754 21248 1792 21282
rect 1826 21248 1832 21282
rect 1714 21209 1832 21248
rect 1714 21175 1720 21209
rect 1754 21175 1792 21209
rect 1826 21175 1832 21209
rect 1714 21136 1832 21175
rect 1714 21102 1720 21136
rect 1754 21102 1792 21136
rect 1826 21102 1832 21136
rect 1714 21070 1832 21102
rect 1594 21043 1640 21055
rect 1714 16472 1832 16473
rect 1202 16466 1832 16472
rect 1202 16432 1244 16466
rect 1278 16432 1320 16466
rect 1354 16432 1395 16466
rect 1429 16432 1470 16466
rect 1504 16432 1545 16466
rect 1579 16432 1620 16466
rect 1654 16432 1695 16466
rect 1729 16432 1832 16466
rect 1090 16417 1832 16432
rect 1090 16394 1792 16417
rect 1090 16360 1168 16394
rect 1202 16360 1246 16394
rect 1280 16360 1324 16394
rect 1358 16360 1402 16394
rect 1436 16360 1480 16394
rect 1514 16360 1558 16394
rect 1592 16360 1636 16394
rect 1670 16360 1714 16394
rect 1748 16383 1792 16394
rect 1826 16383 1832 16417
rect 1748 16360 1832 16383
rect 1090 16354 1832 16360
rect 2020 14640 2072 14646
rect 2020 14565 2072 14588
tri 1984 14490 2020 14526 se
rect 2020 14490 2072 14513
tri 1366 14443 1413 14490 se
rect 1413 14469 2072 14490
rect 1413 14443 2046 14469
tri 2046 14443 2072 14469 nw
rect 2112 14640 2164 14646
rect 2112 14565 2164 14588
tri 1341 14418 1366 14443 se
rect 1366 14438 2041 14443
tri 2041 14438 2046 14443 nw
tri 2107 14438 2112 14443 se
rect 2112 14438 2164 14513
rect 1366 14418 1424 14438
tri 1424 14418 1444 14438 nw
tri 2087 14418 2107 14438 se
rect 2107 14418 2164 14438
rect 1341 14402 1408 14418
tri 1408 14402 1424 14418 nw
tri 2071 14402 2087 14418 se
rect 2087 14402 2164 14418
rect 1341 14302 1393 14402
tri 1393 14387 1408 14402 nw
tri 1490 14387 1505 14402 se
rect 1505 14387 2164 14402
rect 1341 14227 1393 14250
rect 1341 14169 1393 14175
tri 1433 14330 1490 14387 se
rect 1490 14379 2164 14387
rect 1490 14350 2135 14379
tri 2135 14350 2164 14379 nw
rect 1490 14330 1516 14350
tri 1516 14330 1536 14350 nw
rect 1433 14300 1485 14330
tri 1485 14299 1516 14330 nw
rect 1433 14225 1485 14248
rect 1433 14167 1485 14173
rect 507 13226 26404 13232
rect 507 13192 585 13226
rect 619 13192 658 13226
rect 692 13192 731 13226
rect 765 13192 804 13226
rect 507 13154 804 13192
rect 507 9736 513 13154
rect 619 13120 658 13154
rect 692 13120 731 13154
rect 765 13120 804 13154
rect 26326 13154 26404 13226
rect 26326 13120 26364 13154
rect 26398 13120 26404 13154
rect 619 13082 876 13120
rect 691 13048 730 13082
rect 764 13048 803 13082
rect 837 13048 876 13082
rect 26254 13080 26404 13120
rect 26254 13048 26292 13080
rect 691 13046 26292 13048
rect 26326 13046 26364 13080
rect 26398 13046 26404 13080
rect 691 13042 26404 13046
rect 691 9808 697 13042
rect 26214 13008 26404 13042
rect 26214 12974 26220 13008
rect 26254 13006 26404 13008
rect 26254 12974 26292 13006
rect 26214 12972 26292 12974
rect 26326 12972 26364 13006
rect 26398 12972 26404 13006
rect 26214 12934 26404 12972
rect 26214 12900 26220 12934
rect 26254 12932 26404 12934
rect 26254 12900 26292 12932
rect 26214 12898 26292 12900
rect 26326 12898 26364 12932
rect 26398 12898 26404 12932
rect 26214 12860 26404 12898
rect 619 9769 697 9808
rect 619 9736 657 9769
rect 507 9735 657 9736
rect 691 9735 697 9769
rect 507 9697 697 9735
rect 507 9663 513 9697
rect 547 9663 585 9697
rect 619 9696 697 9697
rect 619 9663 657 9696
rect 507 9662 657 9663
rect 691 9662 697 9696
rect 507 9624 697 9662
rect 507 9590 513 9624
rect 547 9590 585 9624
rect 619 9623 697 9624
rect 619 9590 657 9623
rect 507 9589 657 9590
rect 691 9589 697 9623
rect 507 9551 697 9589
rect 507 9517 513 9551
rect 547 9517 585 9551
rect 619 9550 697 9551
rect 619 9517 657 9550
rect 507 9516 657 9517
rect 691 9516 697 9550
rect 507 9478 697 9516
rect 507 9444 513 9478
rect 547 9444 585 9478
rect 619 9477 697 9478
rect 619 9444 657 9477
rect 507 9443 657 9444
rect 691 9443 697 9477
rect 507 9405 697 9443
rect 507 9371 513 9405
rect 547 9371 585 9405
rect 619 9404 697 9405
rect 619 9371 657 9404
rect 507 9370 657 9371
rect 691 9370 697 9404
rect 507 9332 697 9370
rect 507 9298 513 9332
rect 547 9298 585 9332
rect 619 9331 697 9332
rect 619 9298 657 9331
rect 507 9297 657 9298
rect 691 9297 697 9331
rect 507 9259 697 9297
rect 507 9225 513 9259
rect 547 9225 585 9259
rect 619 9258 697 9259
rect 619 9225 657 9258
rect 507 9224 657 9225
rect 691 9224 697 9258
rect 507 9186 697 9224
rect 507 9152 513 9186
rect 547 9152 585 9186
rect 619 9185 697 9186
rect 619 9152 657 9185
rect 507 9151 657 9152
rect 691 9151 697 9185
rect 507 9113 697 9151
rect 507 9079 513 9113
rect 547 9079 585 9113
rect 619 9112 697 9113
rect 619 9079 657 9112
rect 507 9078 657 9079
rect 691 9078 697 9112
rect 507 9040 697 9078
rect 507 9006 513 9040
rect 547 9006 585 9040
rect 619 9039 697 9040
rect 619 9006 657 9039
rect 507 9005 657 9006
rect 691 9005 697 9039
rect 507 8967 697 9005
rect 507 8933 513 8967
rect 547 8933 585 8967
rect 619 8966 697 8967
rect 619 8933 657 8966
rect 507 8932 657 8933
rect 691 8932 697 8966
rect 507 8894 697 8932
rect 507 8860 513 8894
rect 547 8860 585 8894
rect 619 8893 697 8894
rect 619 8860 657 8893
rect 507 8859 657 8860
rect 691 8859 697 8893
rect 507 8821 697 8859
rect 507 8787 513 8821
rect 547 8787 585 8821
rect 619 8820 697 8821
rect 619 8787 657 8820
rect 507 8786 657 8787
rect 691 8786 697 8820
rect 507 8748 697 8786
rect 507 8714 513 8748
rect 547 8714 585 8748
rect 619 8747 697 8748
rect 619 8714 657 8747
rect 507 8713 657 8714
rect 691 8713 697 8747
rect 507 8675 697 8713
rect 507 8641 513 8675
rect 547 8641 585 8675
rect 619 8674 697 8675
rect 619 8641 657 8674
rect 507 8640 657 8641
rect 691 8640 697 8674
rect 507 8602 697 8640
rect 507 8568 513 8602
rect 547 8568 585 8602
rect 619 8601 697 8602
rect 619 8568 657 8601
rect 507 8567 657 8568
rect 691 8567 697 8601
rect 507 8529 697 8567
rect 507 8495 513 8529
rect 547 8495 585 8529
rect 619 8528 697 8529
rect 619 8495 657 8528
rect 507 8494 657 8495
rect 691 8494 697 8528
rect 507 8456 697 8494
rect 507 8422 513 8456
rect 547 8422 585 8456
rect 619 8455 697 8456
rect 619 8422 657 8455
rect 507 8421 657 8422
rect 691 8421 697 8455
rect 507 8383 697 8421
rect 507 8349 513 8383
rect 547 8349 585 8383
rect 619 8382 697 8383
rect 619 8349 657 8382
rect 507 8348 657 8349
rect 691 8348 697 8382
rect 507 8310 697 8348
rect 507 8276 513 8310
rect 547 8276 585 8310
rect 619 8309 697 8310
rect 619 8276 657 8309
rect 507 8275 657 8276
rect 691 8275 697 8309
rect 507 8237 697 8275
rect 507 8203 513 8237
rect 547 8203 585 8237
rect 619 8236 697 8237
rect 619 8203 657 8236
rect 507 8202 657 8203
rect 691 8202 697 8236
rect 507 8164 697 8202
rect 507 8130 513 8164
rect 547 8130 585 8164
rect 619 8163 697 8164
rect 619 8130 657 8163
rect 507 8129 657 8130
rect 691 8129 697 8163
rect 507 8091 697 8129
rect 507 8057 513 8091
rect 547 8057 585 8091
rect 619 8090 697 8091
rect 619 8057 657 8090
rect 507 8056 657 8057
rect 691 8056 697 8090
rect 507 8018 697 8056
rect 507 7984 513 8018
rect 547 7984 585 8018
rect 619 8017 697 8018
rect 619 7984 657 8017
rect 507 7983 657 7984
rect 691 7983 697 8017
rect 507 7945 697 7983
rect 507 7911 513 7945
rect 547 7911 585 7945
rect 619 7944 697 7945
rect 619 7911 657 7944
rect 507 7910 657 7911
rect 691 7910 697 7944
rect 507 7872 697 7910
rect 507 7838 513 7872
rect 547 7838 585 7872
rect 619 7871 697 7872
rect 619 7838 657 7871
rect 507 7837 657 7838
rect 691 7837 697 7871
rect 507 7799 697 7837
rect 507 7765 513 7799
rect 547 7765 585 7799
rect 619 7798 697 7799
rect 619 7765 657 7798
rect 507 7764 657 7765
rect 691 7764 697 7798
rect 507 7726 697 7764
rect 507 7692 513 7726
rect 547 7692 585 7726
rect 619 7725 697 7726
rect 619 7692 657 7725
rect 507 7691 657 7692
rect 691 7691 697 7725
rect 507 7653 697 7691
rect 507 7619 513 7653
rect 547 7619 585 7653
rect 619 7652 697 7653
rect 619 7619 657 7652
rect 507 7618 657 7619
rect 691 7618 697 7652
rect 507 7580 697 7618
rect 507 7546 513 7580
rect 547 7546 585 7580
rect 619 7579 697 7580
rect 619 7546 657 7579
rect 507 7545 657 7546
rect 691 7545 697 7579
rect 507 7507 697 7545
rect 507 7473 513 7507
rect 547 7473 585 7507
rect 619 7506 697 7507
rect 619 7473 657 7506
rect 507 7472 657 7473
rect 691 7472 697 7506
rect 507 7434 697 7472
rect 507 7400 513 7434
rect 547 7400 585 7434
rect 619 7433 697 7434
rect 619 7400 657 7433
rect 507 7399 657 7400
rect 691 7399 697 7433
rect 507 7361 697 7399
rect 507 7327 513 7361
rect 547 7327 585 7361
rect 619 7360 697 7361
rect 619 7327 657 7360
rect 507 7326 657 7327
rect 691 7326 697 7360
rect 507 7288 697 7326
rect 507 7254 513 7288
rect 547 7254 585 7288
rect 619 7287 697 7288
rect 619 7254 657 7287
rect 507 7253 657 7254
rect 691 7253 697 7287
rect 507 7215 697 7253
rect 507 7181 513 7215
rect 547 7181 585 7215
rect 619 7214 697 7215
rect 619 7181 657 7214
rect 507 7180 657 7181
rect 691 7180 697 7214
rect 507 7142 697 7180
rect 507 7108 513 7142
rect 547 7108 585 7142
rect 619 7141 697 7142
rect 619 7108 657 7141
rect 507 7107 657 7108
rect 691 7107 697 7141
rect 507 7069 697 7107
rect 507 7035 513 7069
rect 547 7035 585 7069
rect 619 7068 697 7069
rect 619 7035 657 7068
rect 507 7034 657 7035
rect 691 7034 697 7068
rect 507 6996 697 7034
rect 507 6962 513 6996
rect 547 6962 585 6996
rect 619 6995 697 6996
rect 619 6962 657 6995
rect 507 6961 657 6962
rect 691 6961 697 6995
rect 507 6923 697 6961
rect 507 6889 513 6923
rect 547 6889 585 6923
rect 619 6922 697 6923
rect 619 6889 657 6922
rect 507 6888 657 6889
rect 691 6888 697 6922
rect 507 6850 697 6888
rect 507 6816 513 6850
rect 547 6816 585 6850
rect 619 6849 697 6850
rect 619 6816 657 6849
rect 507 6815 657 6816
rect 691 6815 697 6849
rect 507 6777 697 6815
rect 507 6743 513 6777
rect 547 6743 585 6777
rect 619 6776 697 6777
rect 619 6743 657 6776
rect 507 6742 657 6743
rect 691 6742 697 6776
rect 507 6704 697 6742
rect 507 6670 513 6704
rect 547 6670 585 6704
rect 619 6703 697 6704
rect 619 6670 657 6703
rect 507 6669 657 6670
rect 691 6669 697 6703
rect 507 6631 697 6669
rect 893 12840 26006 12846
rect 893 12806 971 12840
rect 1005 12806 1044 12840
rect 1078 12806 1117 12840
rect 1151 12806 1190 12840
rect 1224 12806 1263 12840
rect 1297 12806 1336 12840
rect 1370 12806 1409 12840
rect 1443 12806 1482 12840
rect 1516 12806 1555 12840
rect 1589 12806 1628 12840
rect 1662 12806 1701 12840
rect 1735 12806 1774 12840
rect 893 12768 1774 12806
rect 893 9638 899 12768
rect 1005 12734 1044 12768
rect 1078 12734 1117 12768
rect 1151 12734 1190 12768
rect 1224 12734 1263 12768
rect 1297 12734 1336 12768
rect 1370 12734 1409 12768
rect 1443 12734 1482 12768
rect 1516 12734 1555 12768
rect 1589 12734 1628 12768
rect 1662 12734 1701 12768
rect 1735 12734 1774 12768
rect 25928 12768 26006 12840
rect 25928 12734 25966 12768
rect 26000 12734 26006 12768
rect 1005 12696 1846 12734
rect 1077 12662 1116 12696
rect 1150 12662 1189 12696
rect 1223 12662 1262 12696
rect 1296 12662 1335 12696
rect 1369 12662 1408 12696
rect 1442 12662 1481 12696
rect 1515 12662 1554 12696
rect 1588 12662 1627 12696
rect 1661 12662 1700 12696
rect 1734 12662 1773 12696
rect 1807 12662 1846 12696
rect 25856 12694 26006 12734
rect 25856 12662 25894 12694
rect 1077 12660 25894 12662
rect 25928 12660 25966 12694
rect 26000 12660 26006 12694
rect 1077 12656 26006 12660
rect 1077 9710 1083 12656
rect 25816 12622 26006 12656
rect 25816 12588 25822 12622
rect 25856 12620 26006 12622
rect 25856 12588 25894 12620
rect 25816 12586 25894 12588
rect 25928 12586 25966 12620
rect 26000 12586 26006 12620
rect 25816 12548 26006 12586
rect 25816 12514 25822 12548
rect 25856 12546 26006 12548
rect 25856 12514 25894 12546
rect 25816 12512 25894 12514
rect 25928 12512 25966 12546
rect 26000 12512 26006 12546
rect 25816 12474 26006 12512
rect 25816 12440 25822 12474
rect 25856 12472 26006 12474
rect 25856 12440 25894 12472
rect 25816 12438 25894 12440
rect 25928 12438 25966 12472
rect 26000 12438 26006 12472
rect 25816 12400 26006 12438
rect 25816 12366 25822 12400
rect 25856 12398 26006 12400
rect 25856 12366 25894 12398
rect 25816 12364 25894 12366
rect 25928 12364 25966 12398
rect 26000 12364 26006 12398
rect 25816 12326 26006 12364
rect 25816 12292 25822 12326
rect 25856 12325 26006 12326
rect 25856 12292 25894 12325
rect 25816 12291 25894 12292
rect 25928 12291 25966 12325
rect 26000 12291 26006 12325
rect 25816 12252 26006 12291
rect 25816 12218 25822 12252
rect 25856 12218 25894 12252
rect 25928 12218 25966 12252
rect 26000 12218 26006 12252
rect 25816 12142 26006 12218
rect 25816 12108 25822 12142
rect 25856 12108 25894 12142
rect 25928 12108 25966 12142
rect 26000 12108 26006 12142
rect 25816 12069 26006 12108
rect 25816 12035 25822 12069
rect 25856 12035 25894 12069
rect 25928 12035 25966 12069
rect 26000 12035 26006 12069
rect 25816 11996 26006 12035
rect 25816 11962 25822 11996
rect 25856 11962 25894 11996
rect 25928 11962 25966 11996
rect 26000 11962 26006 11996
rect 25816 11923 26006 11962
rect 25816 11889 25822 11923
rect 25856 11889 25894 11923
rect 25928 11889 25966 11923
rect 26000 11889 26006 11923
rect 25816 11850 26006 11889
rect 25816 11816 25822 11850
rect 25856 11816 25894 11850
rect 25928 11816 25966 11850
rect 26000 11816 26006 11850
rect 25816 11777 26006 11816
rect 25816 11743 25822 11777
rect 25856 11743 25894 11777
rect 25928 11743 25966 11777
rect 26000 11743 26006 11777
rect 25816 11704 26006 11743
rect 25816 11670 25822 11704
rect 25856 11670 25894 11704
rect 25928 11670 25966 11704
rect 26000 11670 26006 11704
rect 25816 11631 26006 11670
rect 25816 11597 25822 11631
rect 25856 11597 25894 11631
rect 25928 11597 25966 11631
rect 26000 11597 26006 11631
rect 25816 11558 26006 11597
rect 25816 11524 25822 11558
rect 25856 11524 25894 11558
rect 25928 11524 25966 11558
rect 26000 11524 26006 11558
rect 25816 11485 26006 11524
rect 25816 11451 25822 11485
rect 25856 11451 25894 11485
rect 25928 11451 25966 11485
rect 26000 11451 26006 11485
rect 25816 11412 26006 11451
rect 25816 11378 25822 11412
rect 25856 11378 25894 11412
rect 25928 11378 25966 11412
rect 26000 11378 26006 11412
rect 25816 11339 26006 11378
rect 25816 11305 25822 11339
rect 25856 11305 25894 11339
rect 25928 11305 25966 11339
rect 26000 11305 26006 11339
rect 25816 11266 26006 11305
rect 25816 11232 25822 11266
rect 25856 11232 25894 11266
rect 25928 11232 25966 11266
rect 26000 11232 26006 11266
rect 25816 11193 26006 11232
rect 25816 11159 25822 11193
rect 25856 11159 25894 11193
rect 25928 11159 25966 11193
rect 26000 11159 26006 11193
rect 25816 11120 26006 11159
rect 25816 11086 25822 11120
rect 25856 11086 25894 11120
rect 25928 11086 25966 11120
rect 26000 11086 26006 11120
rect 25816 11047 26006 11086
rect 25816 11013 25822 11047
rect 25856 11013 25894 11047
rect 25928 11013 25966 11047
rect 26000 11013 26006 11047
rect 25816 10974 26006 11013
rect 25816 10940 25822 10974
rect 25856 10940 25894 10974
rect 25928 10940 25966 10974
rect 26000 10940 26006 10974
rect 25816 10901 26006 10940
rect 25816 10867 25822 10901
rect 25856 10867 25894 10901
rect 25928 10867 25966 10901
rect 26000 10867 26006 10901
rect 25816 10828 26006 10867
rect 25816 10794 25822 10828
rect 25856 10794 25894 10828
rect 25928 10794 25966 10828
rect 26000 10794 26006 10828
rect 1341 10756 1730 10762
rect 1393 10704 1678 10756
rect 1341 10689 1409 10704
rect 1393 10682 1409 10689
tri 1409 10682 1431 10704 nw
tri 1632 10682 1654 10704 ne
rect 1654 10689 1730 10704
rect 1654 10682 1678 10689
tri 1393 10666 1409 10682 nw
tri 1654 10666 1670 10682 ne
rect 1670 10666 1678 10682
tri 1670 10658 1678 10666 ne
rect 1341 10631 1393 10637
rect 1678 10631 1730 10637
rect 25816 10755 26006 10794
rect 25816 10721 25822 10755
rect 25856 10721 25894 10755
rect 25928 10721 25966 10755
rect 26000 10721 26006 10755
rect 25816 10682 26006 10721
rect 25816 10648 25822 10682
rect 25856 10648 25894 10682
rect 25928 10648 25966 10682
rect 26000 10648 26006 10682
rect 25816 10609 26006 10648
rect 1289 10584 2086 10590
rect 1289 10550 1301 10584
rect 1335 10550 1382 10584
rect 1416 10550 1462 10584
rect 1496 10550 1542 10584
rect 1576 10550 1622 10584
rect 1656 10550 1702 10584
rect 1736 10550 1782 10584
rect 1816 10550 1862 10584
rect 1896 10550 1942 10584
rect 1976 10575 2086 10584
tri 2086 10575 2101 10590 sw
rect 25816 10575 25822 10609
rect 25856 10575 25894 10609
rect 25928 10575 25966 10609
rect 26000 10575 26006 10609
rect 1976 10550 2101 10575
rect 1289 10547 2101 10550
tri 2101 10547 2129 10575 sw
rect 1289 10544 2471 10547
tri 2050 10536 2058 10544 ne
rect 2058 10541 2471 10544
rect 2058 10536 2419 10541
tri 2058 10511 2083 10536 ne
rect 2083 10511 2419 10536
rect 1678 10505 2039 10511
tri 2083 10509 2085 10511 ne
rect 2085 10509 2419 10511
rect 1730 10499 2039 10505
rect 1730 10465 1999 10499
rect 2033 10465 2039 10499
rect 1730 10453 2039 10465
rect 1678 10435 2039 10453
rect 1730 10426 2039 10435
rect 1730 10392 1999 10426
rect 2033 10392 2039 10426
rect 2419 10477 2471 10489
rect 2419 10419 2471 10425
rect 25816 10536 26006 10575
rect 25816 10502 25822 10536
rect 25856 10502 25894 10536
rect 25928 10502 25966 10536
rect 26000 10502 26006 10536
rect 25816 10463 26006 10502
rect 25816 10429 25822 10463
rect 25856 10429 25894 10463
rect 25928 10429 25966 10463
rect 26000 10429 26006 10463
rect 1730 10383 2039 10392
rect 1678 10364 2039 10383
rect 1730 10352 2039 10364
rect 1730 10318 1999 10352
rect 2033 10318 2039 10352
rect 1730 10312 2039 10318
rect 1678 10306 2039 10312
rect 25816 10390 26006 10429
rect 25816 10356 25822 10390
rect 25856 10356 25894 10390
rect 25928 10356 25966 10390
rect 26000 10356 26006 10390
rect 25816 10317 26006 10356
rect 25816 10283 25822 10317
rect 25856 10283 25894 10317
rect 25928 10283 25966 10317
rect 26000 10283 26006 10317
rect 25816 10244 26006 10283
rect 25816 10210 25822 10244
rect 25856 10210 25894 10244
rect 25928 10210 25966 10244
rect 26000 10210 26006 10244
rect 25816 10171 26006 10210
rect 1837 10149 1883 10161
rect 1837 10115 1843 10149
rect 1877 10115 1883 10149
rect 1837 10080 1883 10115
rect 25816 10137 25822 10171
rect 25856 10137 25894 10171
rect 25928 10137 25966 10171
rect 26000 10137 26006 10171
rect 25816 10098 26006 10137
rect 1163 10077 2223 10080
rect 1163 10074 1843 10077
rect 1215 10043 1843 10074
rect 1877 10074 2223 10077
rect 1877 10043 2171 10074
rect 1215 10030 2171 10043
rect 1163 10010 1215 10022
rect 1163 9952 1215 9958
rect 2171 10010 2223 10022
rect 2171 9952 2223 9958
rect 25816 10064 25822 10098
rect 25856 10064 25894 10098
rect 25928 10064 25966 10098
rect 26000 10064 26006 10098
rect 25816 10025 26006 10064
rect 25816 9991 25822 10025
rect 25856 9991 25894 10025
rect 25928 9991 25966 10025
rect 26000 9991 26006 10025
rect 25816 9952 26006 9991
rect 25816 9918 25822 9952
rect 25856 9918 25894 9952
rect 25928 9918 25966 9952
rect 26000 9918 26006 9952
rect 25816 9879 26006 9918
rect 2419 9870 2471 9876
rect 2419 9806 2471 9818
rect 1289 9788 2419 9794
rect 1289 9754 1301 9788
rect 1335 9754 1400 9788
rect 1434 9754 1499 9788
rect 1533 9754 2419 9788
rect 1289 9748 2471 9754
rect 25816 9845 25822 9879
rect 25856 9845 25894 9879
rect 25928 9845 25966 9879
rect 26000 9845 26006 9879
rect 25816 9806 26006 9845
rect 25816 9772 25822 9806
rect 25856 9772 25894 9806
rect 25928 9772 25966 9806
rect 26000 9772 26006 9806
rect 1005 9671 1083 9710
rect 25816 9733 26006 9772
rect 1005 9638 1043 9671
rect 893 9637 1043 9638
rect 1077 9637 1083 9671
rect 893 9599 1083 9637
rect 893 9565 899 9599
rect 933 9565 971 9599
rect 1005 9598 1083 9599
rect 1005 9565 1043 9598
rect 893 9564 1043 9565
rect 1077 9564 1083 9598
rect 893 9526 1083 9564
rect 893 9492 899 9526
rect 933 9492 971 9526
rect 1005 9525 1083 9526
rect 1005 9492 1043 9525
rect 893 9491 1043 9492
rect 1077 9491 1083 9525
rect 1238 9697 1596 9703
rect 1238 9691 1433 9697
rect 1238 9657 1244 9691
rect 1278 9657 1433 9691
rect 1238 9645 1433 9657
rect 1485 9691 1596 9697
rect 1485 9657 1556 9691
rect 1590 9657 1596 9691
rect 1485 9645 1596 9657
rect 1238 9627 1596 9645
rect 1238 9618 1433 9627
rect 1238 9584 1244 9618
rect 1278 9584 1433 9618
rect 1238 9575 1433 9584
rect 1485 9618 1596 9627
rect 1485 9584 1556 9618
rect 1590 9584 1596 9618
rect 1485 9575 1596 9584
rect 1238 9556 1596 9575
rect 1238 9544 1433 9556
rect 1238 9510 1244 9544
rect 1278 9510 1433 9544
rect 1238 9504 1433 9510
rect 1485 9544 1596 9556
rect 1485 9510 1556 9544
rect 1590 9510 1596 9544
rect 25816 9699 25822 9733
rect 25856 9699 25894 9733
rect 25928 9699 25966 9733
rect 26000 9699 26006 9733
rect 25816 9660 26006 9699
rect 25816 9626 25822 9660
rect 25856 9626 25894 9660
rect 25928 9626 25966 9660
rect 26000 9626 26006 9660
rect 25816 9587 26006 9626
rect 25816 9553 25822 9587
rect 25856 9553 25894 9587
rect 25928 9553 25966 9587
rect 26000 9553 26006 9587
rect 1485 9504 1596 9510
rect 1238 9498 1596 9504
rect 2337 9514 2389 9520
rect 893 9453 1083 9491
rect 893 9419 899 9453
rect 933 9419 971 9453
rect 1005 9452 1083 9453
rect 1005 9419 1043 9452
rect 893 9418 1043 9419
rect 1077 9418 1083 9452
rect 893 9380 1083 9418
rect 893 9346 899 9380
rect 933 9346 971 9380
rect 1005 9379 1083 9380
rect 1005 9346 1043 9379
rect 893 9345 1043 9346
rect 1077 9345 1083 9379
rect 893 9307 1083 9345
rect 1163 9462 2337 9466
rect 1163 9460 2389 9462
rect 1215 9454 2389 9460
rect 1215 9420 1400 9454
rect 1434 9450 2389 9454
rect 1434 9420 2337 9450
rect 1215 9416 2337 9420
rect 1163 9396 1215 9408
rect 1163 9338 1215 9344
rect 1394 9382 1440 9416
rect 2337 9392 2389 9398
rect 25816 9514 26006 9553
rect 25816 9480 25822 9514
rect 25856 9480 25894 9514
rect 25928 9480 25966 9514
rect 26000 9480 26006 9514
rect 25816 9441 26006 9480
rect 25816 9407 25822 9441
rect 25856 9407 25894 9441
rect 25928 9407 25966 9441
rect 26000 9407 26006 9441
rect 1394 9348 1400 9382
rect 1434 9348 1440 9382
rect 1394 9336 1440 9348
rect 25816 9368 26006 9407
rect 893 9273 899 9307
rect 933 9273 971 9307
rect 1005 9306 1083 9307
rect 1005 9273 1043 9306
rect 893 9272 1043 9273
rect 1077 9272 1083 9306
rect 893 9234 1083 9272
rect 893 9200 899 9234
rect 933 9200 971 9234
rect 1005 9233 1083 9234
rect 1005 9200 1043 9233
rect 893 9199 1043 9200
rect 1077 9199 1083 9233
rect 893 9161 1083 9199
rect 893 9127 899 9161
rect 933 9127 971 9161
rect 1005 9160 1083 9161
rect 1005 9127 1043 9160
rect 893 9126 1043 9127
rect 1077 9126 1083 9160
rect 893 9088 1083 9126
rect 893 9054 899 9088
rect 933 9054 971 9088
rect 1005 9087 1083 9088
rect 1005 9054 1043 9087
rect 893 9053 1043 9054
rect 1077 9053 1083 9087
rect 893 9015 1083 9053
rect 893 8981 899 9015
rect 933 8981 971 9015
rect 1005 9014 1083 9015
rect 1005 8981 1043 9014
rect 893 8980 1043 8981
rect 1077 8980 1083 9014
rect 893 8942 1083 8980
rect 893 8908 899 8942
rect 933 8908 971 8942
rect 1005 8941 1083 8942
rect 1005 8908 1043 8941
rect 893 8907 1043 8908
rect 1077 8907 1083 8941
rect 893 8869 1083 8907
rect 893 8835 899 8869
rect 933 8835 971 8869
rect 1005 8868 1083 8869
rect 1005 8835 1043 8868
rect 893 8834 1043 8835
rect 1077 8834 1083 8868
rect 893 8796 1083 8834
rect 893 8762 899 8796
rect 933 8762 971 8796
rect 1005 8795 1083 8796
rect 1005 8762 1043 8795
rect 893 8761 1043 8762
rect 1077 8761 1083 8795
rect 893 8723 1083 8761
rect 893 8689 899 8723
rect 933 8689 971 8723
rect 1005 8722 1083 8723
rect 1005 8689 1043 8722
rect 893 8688 1043 8689
rect 1077 8688 1083 8722
rect 893 8650 1083 8688
rect 893 8616 899 8650
rect 933 8616 971 8650
rect 1005 8649 1083 8650
rect 1005 8616 1043 8649
rect 893 8615 1043 8616
rect 1077 8615 1083 8649
rect 893 8577 1083 8615
rect 893 8543 899 8577
rect 933 8543 971 8577
rect 1005 8576 1083 8577
rect 1005 8543 1043 8576
rect 893 8542 1043 8543
rect 1077 8542 1083 8576
rect 893 8504 1083 8542
rect 893 8470 899 8504
rect 933 8470 971 8504
rect 1005 8503 1083 8504
rect 1005 8470 1043 8503
rect 893 8469 1043 8470
rect 1077 8469 1083 8503
rect 893 8431 1083 8469
rect 893 8397 899 8431
rect 933 8397 971 8431
rect 1005 8430 1083 8431
rect 1005 8397 1043 8430
rect 893 8396 1043 8397
rect 1077 8396 1083 8430
rect 893 8358 1083 8396
rect 893 8324 899 8358
rect 933 8324 971 8358
rect 1005 8357 1083 8358
rect 1005 8324 1043 8357
rect 893 8323 1043 8324
rect 1077 8323 1083 8357
rect 893 8285 1083 8323
rect 893 8251 899 8285
rect 933 8251 971 8285
rect 1005 8284 1083 8285
rect 1005 8251 1043 8284
rect 893 8250 1043 8251
rect 1077 8250 1083 8284
rect 893 8212 1083 8250
rect 893 8178 899 8212
rect 933 8178 971 8212
rect 1005 8211 1083 8212
rect 1005 8178 1043 8211
rect 893 8177 1043 8178
rect 1077 8177 1083 8211
rect 893 8139 1083 8177
rect 893 8105 899 8139
rect 933 8105 971 8139
rect 1005 8138 1083 8139
rect 1005 8105 1043 8138
rect 893 8104 1043 8105
rect 1077 8104 1083 8138
rect 893 8066 1083 8104
rect 893 8032 899 8066
rect 933 8032 971 8066
rect 1005 8065 1083 8066
rect 1005 8032 1043 8065
rect 893 8031 1043 8032
rect 1077 8031 1083 8065
rect 893 7993 1083 8031
rect 893 7959 899 7993
rect 933 7959 971 7993
rect 1005 7992 1083 7993
rect 1005 7959 1043 7992
rect 893 7958 1043 7959
rect 1077 7958 1083 7992
rect 893 7920 1083 7958
rect 893 7886 899 7920
rect 933 7886 971 7920
rect 1005 7919 1083 7920
rect 1005 7886 1043 7919
rect 893 7885 1043 7886
rect 1077 7885 1083 7919
rect 25816 9334 25822 9368
rect 25856 9334 25894 9368
rect 25928 9334 25966 9368
rect 26000 9334 26006 9368
rect 25816 9295 26006 9334
rect 25816 9261 25822 9295
rect 25856 9261 25894 9295
rect 25928 9261 25966 9295
rect 26000 9261 26006 9295
rect 25816 9222 26006 9261
rect 25816 9188 25822 9222
rect 25856 9188 25894 9222
rect 25928 9188 25966 9222
rect 26000 9188 26006 9222
rect 25816 9149 26006 9188
rect 25816 9115 25822 9149
rect 25856 9115 25894 9149
rect 25928 9115 25966 9149
rect 26000 9115 26006 9149
rect 25816 9076 26006 9115
rect 25816 9042 25822 9076
rect 25856 9042 25894 9076
rect 25928 9042 25966 9076
rect 26000 9042 26006 9076
rect 25816 9003 26006 9042
rect 25816 8969 25822 9003
rect 25856 8969 25894 9003
rect 25928 8969 25966 9003
rect 26000 8969 26006 9003
rect 25816 8930 26006 8969
rect 25816 8896 25822 8930
rect 25856 8896 25894 8930
rect 25928 8896 25966 8930
rect 26000 8896 26006 8930
rect 25816 8857 26006 8896
rect 25816 8823 25822 8857
rect 25856 8823 25894 8857
rect 25928 8823 25966 8857
rect 26000 8823 26006 8857
rect 25816 8784 26006 8823
rect 25816 8750 25822 8784
rect 25856 8750 25894 8784
rect 25928 8750 25966 8784
rect 26000 8750 26006 8784
rect 25816 8711 26006 8750
rect 25816 8677 25822 8711
rect 25856 8677 25894 8711
rect 25928 8677 25966 8711
rect 26000 8677 26006 8711
rect 25816 8638 26006 8677
rect 25816 8604 25822 8638
rect 25856 8604 25894 8638
rect 25928 8604 25966 8638
rect 26000 8604 26006 8638
rect 25816 8565 26006 8604
rect 25816 8531 25822 8565
rect 25856 8531 25894 8565
rect 25928 8531 25966 8565
rect 26000 8531 26006 8565
rect 25816 8492 26006 8531
rect 25816 8458 25822 8492
rect 25856 8458 25894 8492
rect 25928 8458 25966 8492
rect 26000 8458 26006 8492
rect 25816 8419 26006 8458
rect 25816 8385 25822 8419
rect 25856 8385 25894 8419
rect 25928 8385 25966 8419
rect 26000 8385 26006 8419
rect 25816 8346 26006 8385
rect 25816 8312 25822 8346
rect 25856 8312 25894 8346
rect 25928 8312 25966 8346
rect 26000 8312 26006 8346
rect 25816 8273 26006 8312
rect 25816 8239 25822 8273
rect 25856 8239 25894 8273
rect 25928 8239 25966 8273
rect 26000 8239 26006 8273
rect 25816 8200 26006 8239
rect 25816 8166 25822 8200
rect 25856 8166 25894 8200
rect 25928 8166 25966 8200
rect 26000 8166 26006 8200
rect 25816 8127 26006 8166
rect 25816 8093 25822 8127
rect 25856 8093 25894 8127
rect 25928 8093 25966 8127
rect 26000 8093 26006 8127
rect 25816 8054 26006 8093
rect 25816 8020 25822 8054
rect 25856 8020 25894 8054
rect 25928 8020 25966 8054
rect 26000 8020 26006 8054
rect 25816 7981 26006 8020
rect 25816 7947 25822 7981
rect 25856 7947 25894 7981
rect 25928 7947 25966 7981
rect 26000 7947 26006 7981
rect 25816 7908 26006 7947
rect 893 7847 1083 7885
rect 893 7813 899 7847
rect 933 7813 971 7847
rect 1005 7846 1083 7847
rect 1005 7813 1043 7846
rect 893 7812 1043 7813
rect 1077 7812 1083 7846
tri 7981 7883 7984 7886 se
rect 7984 7883 8656 7886
tri 8656 7883 8659 7886 sw
rect 7981 7837 8659 7883
tri 7981 7835 7983 7837 ne
rect 7983 7835 8657 7837
tri 8657 7835 8659 7837 nw
tri 9485 7883 9488 7886 se
rect 9488 7883 9903 7886
tri 9903 7883 9906 7886 sw
tri 12958 7883 12961 7886 se
rect 12961 7883 13376 7886
tri 13376 7883 13379 7886 sw
rect 9485 7837 9906 7883
rect 11286 7837 11593 7883
rect 12958 7837 13379 7883
tri 9485 7835 9487 7837 ne
rect 9487 7835 9904 7837
tri 9904 7835 9906 7837 nw
tri 12958 7835 12960 7837 ne
rect 12960 7835 13377 7837
tri 13377 7835 13379 7837 nw
tri 14205 7883 14208 7886 se
rect 14208 7883 14880 7886
tri 14880 7883 14883 7886 sw
rect 14205 7837 14883 7883
tri 14205 7835 14207 7837 ne
rect 14207 7835 14881 7837
tri 14881 7835 14883 7837 nw
rect 25816 7874 25822 7908
rect 25856 7874 25894 7908
rect 25928 7874 25966 7908
rect 26000 7874 26006 7908
rect 25816 7835 26006 7874
tri 7983 7834 7984 7835 ne
rect 7984 7834 8656 7835
tri 8656 7834 8657 7835 nw
tri 9487 7834 9488 7835 ne
rect 9488 7834 9903 7835
tri 9903 7834 9904 7835 nw
tri 12960 7834 12961 7835 ne
rect 12961 7834 13376 7835
tri 13376 7834 13377 7835 nw
tri 14207 7834 14208 7835 ne
rect 14208 7834 14880 7835
tri 14880 7834 14881 7835 nw
rect 893 7774 1083 7812
rect 893 7740 899 7774
rect 933 7740 971 7774
rect 1005 7773 1083 7774
rect 1005 7740 1043 7773
rect 893 7739 1043 7740
rect 1077 7739 1083 7773
rect 893 7701 1083 7739
rect 893 7667 899 7701
rect 933 7667 971 7701
rect 1005 7700 1083 7701
rect 1005 7667 1043 7700
rect 893 7666 1043 7667
rect 1077 7666 1083 7700
rect 893 7628 1083 7666
rect 893 7594 899 7628
rect 933 7594 971 7628
rect 1005 7627 1083 7628
rect 1005 7594 1043 7627
rect 893 7593 1043 7594
rect 1077 7593 1083 7627
rect 893 7555 1083 7593
rect 893 7521 899 7555
rect 933 7521 971 7555
rect 1005 7554 1083 7555
rect 1005 7521 1043 7554
rect 893 7520 1043 7521
rect 1077 7520 1083 7554
rect 893 7482 1083 7520
rect 893 7448 899 7482
rect 933 7448 971 7482
rect 1005 7481 1083 7482
rect 1005 7448 1043 7481
rect 893 7447 1043 7448
rect 1077 7447 1083 7481
rect 893 7409 1083 7447
rect 893 7375 899 7409
rect 933 7375 971 7409
rect 1005 7408 1083 7409
rect 1005 7375 1043 7408
rect 893 7374 1043 7375
rect 1077 7374 1083 7408
rect 893 7336 1083 7374
rect 893 7302 899 7336
rect 933 7302 971 7336
rect 1005 7335 1083 7336
rect 1005 7302 1043 7335
rect 893 7301 1043 7302
rect 1077 7301 1083 7335
rect 893 7263 1083 7301
rect 893 7229 899 7263
rect 933 7229 971 7263
rect 1005 7262 1083 7263
rect 1005 7229 1043 7262
rect 893 7228 1043 7229
rect 1077 7228 1083 7262
rect 893 7190 1083 7228
rect 893 7156 899 7190
rect 933 7156 971 7190
rect 1005 7189 1083 7190
rect 1005 7156 1043 7189
rect 893 7155 1043 7156
rect 1077 7155 1083 7189
rect 893 7117 1083 7155
rect 893 7083 899 7117
rect 933 7083 971 7117
rect 1005 7116 1083 7117
rect 1005 7083 1043 7116
rect 893 7082 1043 7083
rect 1077 7082 1083 7116
rect 893 7044 1083 7082
rect 893 7010 899 7044
rect 933 7010 971 7044
rect 1005 7043 1083 7044
rect 1005 7010 1043 7043
rect 893 7009 1043 7010
rect 1077 7009 1083 7043
rect 893 6971 1083 7009
rect 893 6937 899 6971
rect 933 6937 971 6971
rect 1005 6970 1083 6971
rect 1005 6937 1043 6970
rect 893 6936 1043 6937
rect 1077 6936 1083 6970
rect 893 6898 1083 6936
rect 893 6864 899 6898
rect 933 6864 971 6898
rect 1005 6897 1083 6898
rect 1005 6864 1043 6897
rect 893 6863 1043 6864
rect 1077 6863 1083 6897
rect 893 6830 1083 6863
rect 25816 7801 25822 7835
rect 25856 7801 25894 7835
rect 25928 7801 25966 7835
rect 26000 7801 26006 7835
rect 25816 7762 26006 7801
rect 25816 7728 25822 7762
rect 25856 7728 25894 7762
rect 25928 7728 25966 7762
rect 26000 7728 26006 7762
rect 25816 7689 26006 7728
rect 25816 7655 25822 7689
rect 25856 7655 25894 7689
rect 25928 7655 25966 7689
rect 26000 7655 26006 7689
rect 25816 7616 26006 7655
rect 25816 6830 25822 7616
rect 893 6825 25822 6830
rect 893 6791 899 6825
rect 933 6791 971 6825
rect 1005 6824 25822 6825
rect 1005 6791 1043 6824
rect 893 6752 1043 6791
rect 25053 6790 25092 6824
rect 25126 6790 25165 6824
rect 25199 6790 25238 6824
rect 25272 6790 25311 6824
rect 25345 6790 25384 6824
rect 25418 6790 25457 6824
rect 25491 6790 25530 6824
rect 25564 6790 25603 6824
rect 25637 6790 25676 6824
rect 25710 6790 25749 6824
rect 25783 6790 25822 6824
rect 25053 6752 25894 6790
rect 893 6718 899 6752
rect 933 6718 971 6752
rect 893 6646 971 6718
rect 25125 6718 25164 6752
rect 25198 6718 25237 6752
rect 25271 6718 25310 6752
rect 25344 6718 25383 6752
rect 25417 6718 25456 6752
rect 25490 6718 25529 6752
rect 25563 6718 25602 6752
rect 25636 6718 25675 6752
rect 25709 6718 25748 6752
rect 25782 6718 25821 6752
rect 25855 6718 25894 6752
rect 26000 6718 26006 7616
rect 25125 6680 26006 6718
rect 25125 6646 25164 6680
rect 25198 6646 25237 6680
rect 25271 6646 25310 6680
rect 25344 6646 25383 6680
rect 25417 6646 25456 6680
rect 25490 6646 25529 6680
rect 25563 6646 25602 6680
rect 25636 6646 25675 6680
rect 25709 6646 25748 6680
rect 25782 6646 25821 6680
rect 25855 6646 25894 6680
rect 25928 6646 26006 6680
rect 893 6640 26006 6646
rect 26214 12826 26220 12860
rect 26254 12858 26404 12860
rect 26254 12826 26292 12858
rect 26214 12824 26292 12826
rect 26326 12824 26364 12858
rect 26398 12824 26404 12858
rect 26214 12786 26404 12824
rect 26214 12752 26220 12786
rect 26254 12784 26404 12786
rect 26254 12752 26292 12784
rect 26214 12750 26292 12752
rect 26326 12750 26364 12784
rect 26398 12750 26404 12784
rect 26214 12712 26404 12750
rect 26214 12678 26220 12712
rect 26254 12711 26404 12712
rect 26254 12678 26292 12711
rect 26214 12677 26292 12678
rect 26326 12677 26364 12711
rect 26398 12677 26404 12711
rect 26214 12638 26404 12677
rect 26214 12604 26220 12638
rect 26254 12604 26292 12638
rect 26326 12604 26364 12638
rect 26398 12604 26404 12638
rect 26214 12528 26404 12604
rect 26214 12494 26220 12528
rect 26254 12494 26292 12528
rect 26326 12494 26364 12528
rect 26398 12494 26404 12528
rect 26214 12455 26404 12494
rect 26214 12421 26220 12455
rect 26254 12421 26292 12455
rect 26326 12421 26364 12455
rect 26398 12421 26404 12455
rect 26214 12382 26404 12421
rect 26214 12348 26220 12382
rect 26254 12348 26292 12382
rect 26326 12348 26364 12382
rect 26398 12348 26404 12382
rect 26214 12309 26404 12348
rect 26214 12275 26220 12309
rect 26254 12275 26292 12309
rect 26326 12275 26364 12309
rect 26398 12275 26404 12309
rect 26214 12236 26404 12275
rect 26214 12202 26220 12236
rect 26254 12202 26292 12236
rect 26326 12202 26364 12236
rect 26398 12202 26404 12236
rect 26214 12163 26404 12202
rect 507 6597 513 6631
rect 547 6597 585 6631
rect 619 6630 697 6631
rect 619 6597 657 6630
rect 507 6596 657 6597
rect 691 6596 697 6630
rect 507 6558 697 6596
rect 507 6524 513 6558
rect 547 6524 585 6558
rect 619 6557 697 6558
rect 619 6524 657 6557
rect 507 6523 657 6524
rect 691 6523 697 6557
rect 507 6485 697 6523
rect 507 6451 513 6485
rect 547 6451 585 6485
rect 619 6484 697 6485
rect 619 6451 657 6484
rect 507 6450 657 6451
rect 691 6450 697 6484
rect 507 6412 697 6450
rect 507 6378 513 6412
rect 547 6378 585 6412
rect 619 6411 697 6412
rect 619 6378 657 6411
rect 507 6377 657 6378
rect 691 6377 697 6411
rect 507 6339 697 6377
rect 507 6305 513 6339
rect 547 6305 585 6339
rect 619 6338 697 6339
rect 619 6305 657 6338
rect 507 6304 657 6305
rect 691 6304 697 6338
tri 24932 6333 24987 6388 se
rect 24987 6336 25526 6388
rect 25578 6336 25590 6388
rect 25642 6336 25648 6388
rect 24987 6333 25005 6336
tri 25005 6333 25008 6336 nw
rect 507 6266 697 6304
rect 2094 6281 2100 6333
rect 2152 6281 2164 6333
rect 2216 6303 24975 6333
tri 24975 6303 25005 6333 nw
rect 2216 6281 2222 6303
rect 25063 6275 25069 6293
rect 507 6232 513 6266
rect 547 6232 585 6266
rect 619 6265 697 6266
rect 619 6232 657 6265
rect 507 6231 657 6232
rect 691 6231 697 6265
rect 507 6193 697 6231
rect 1926 6207 1932 6259
rect 1984 6207 1996 6259
rect 2048 6241 2054 6259
rect 2295 6241 25069 6275
rect 25121 6241 25133 6293
rect 25185 6241 25191 6293
rect 2048 6207 2329 6241
rect 507 6159 513 6193
rect 547 6159 585 6193
rect 619 6192 697 6193
rect 619 6159 657 6192
rect 507 6158 657 6159
rect 691 6158 697 6192
rect 507 6120 697 6158
rect 507 6086 513 6120
rect 547 6086 585 6120
rect 619 6119 697 6120
rect 619 6086 657 6119
rect 507 6085 657 6086
rect 691 6085 697 6119
rect 507 6047 697 6085
rect 507 6013 513 6047
rect 547 6013 585 6047
rect 619 6046 697 6047
rect 619 6013 657 6046
rect 507 6012 657 6013
rect 691 6012 697 6046
rect 507 5974 697 6012
rect 507 5940 513 5974
rect 547 5940 585 5974
rect 619 5973 697 5974
rect 619 5940 657 5973
rect 507 5939 657 5940
rect 691 5939 697 5973
rect 507 5901 697 5939
rect 507 5867 513 5901
rect 547 5867 585 5901
rect 619 5900 697 5901
rect 619 5867 657 5900
rect 507 5866 657 5867
rect 691 5866 697 5900
rect 2255 5993 2307 5994
rect 2255 5988 8667 5993
rect 2307 5948 8667 5988
rect 2255 5924 2307 5936
tri 2307 5922 2333 5948 nw
rect 8661 5941 8667 5948
rect 8719 5941 8731 5993
rect 8783 5941 8789 5993
rect 2255 5866 2307 5872
rect 2353 5866 2359 5918
rect 2411 5866 2423 5918
rect 2475 5910 8607 5918
tri 8607 5910 8615 5918 sw
tri 8805 5910 8813 5918 se
rect 8813 5910 13064 5918
rect 2475 5866 13064 5910
rect 13116 5866 13128 5918
rect 13180 5866 13186 5918
rect 507 5833 697 5866
rect 26214 5833 26220 12163
rect 507 5828 26220 5833
rect 507 5794 513 5828
rect 547 5794 585 5828
rect 619 5827 26220 5828
rect 619 5794 657 5827
rect 507 5755 657 5794
rect 26035 5793 26074 5827
rect 26108 5793 26147 5827
rect 26181 5793 26220 5827
rect 26035 5755 26292 5793
rect 507 5721 513 5755
rect 547 5721 585 5755
rect 507 5649 585 5721
rect 26107 5721 26146 5755
rect 26180 5721 26219 5755
rect 26253 5721 26292 5755
rect 26398 5721 26404 12163
rect 26107 5683 26404 5721
rect 26107 5649 26146 5683
rect 26180 5649 26219 5683
rect 26253 5649 26292 5683
rect 26326 5649 26404 5683
rect 507 5643 26404 5649
rect 7882 5236 25468 5242
rect 7882 5210 25416 5236
rect 7882 5201 8010 5210
tri 7321 5182 7340 5201 se
rect 7340 5182 7348 5201
tri 7289 5150 7321 5182 se
rect 7321 5150 7348 5182
tri 7248 5109 7289 5150 se
rect 7289 5149 7348 5150
rect 7400 5149 7412 5201
rect 7464 5149 7470 5201
rect 7882 5149 7888 5201
rect 7940 5149 7952 5201
rect 8004 5149 8010 5201
rect 12321 5176 25377 5182
rect 12321 5150 25325 5176
rect 7289 5148 7470 5149
rect 7289 5109 7467 5148
tri 7467 5145 7470 5148 nw
rect 12321 5109 12384 5150
rect 25325 5096 25377 5124
rect 25416 5156 25468 5184
rect 25416 5098 25468 5104
rect 25325 5038 25377 5044
rect 118 4217 523 4707
rect 24702 4136 24991 4263
rect 7531 3728 7598 3930
rect 8440 3606 17159 3682
rect 2255 3501 2320 3552
rect -968 3040 -962 3092
rect -910 3040 -877 3092
rect -825 3040 -819 3092
rect -968 3012 -819 3040
rect -968 2960 -962 3012
rect -910 2960 -877 3012
rect -825 2960 -819 3012
rect -968 2932 -819 2960
rect -631 3066 -231 3072
rect -631 3032 -619 3066
rect -585 3056 -533 3066
rect -499 3056 -447 3066
rect -413 3056 -362 3066
rect -328 3056 -277 3066
rect -243 3056 -231 3066
rect -631 3004 -617 3032
rect -565 3004 -535 3056
rect -483 3004 -453 3056
rect -401 3004 -371 3056
rect -319 3004 -289 3056
rect -237 3004 -231 3056
rect -631 2988 -231 3004
rect -631 2954 -619 2988
rect -585 2954 -533 2988
rect -499 2954 -447 2988
rect -413 2954 -362 2988
rect -328 2954 -277 2988
rect -243 2954 -231 2988
rect -631 2948 -231 2954
rect -151 3066 249 3072
rect -151 3037 -139 3066
rect -105 3037 -53 3066
rect -19 3037 33 3066
rect 67 3037 118 3066
rect -151 2985 -141 3037
rect -89 2985 -65 3037
rect -13 2985 11 3037
rect 67 3032 86 3037
rect 152 3032 203 3066
rect 237 3032 249 3066
rect 63 2988 86 3032
rect 138 2988 249 3032
rect 67 2985 86 2988
rect -151 2954 -139 2985
rect -105 2954 -53 2985
rect -19 2954 33 2985
rect 67 2954 118 2985
rect 152 2954 203 2988
rect 237 2954 249 2988
rect -151 2948 249 2954
rect 334 3066 734 3072
rect 334 3032 346 3066
rect 380 3037 432 3066
rect 466 3037 518 3066
rect 552 3037 603 3066
rect 409 3032 432 3037
rect 334 2988 357 3032
rect 409 2988 433 3032
rect 334 2954 346 2988
rect 409 2985 432 2988
rect 485 2985 509 3037
rect 561 2985 584 3037
rect 637 3032 688 3066
rect 722 3032 734 3066
rect 636 2988 734 3032
rect 380 2954 432 2985
rect 466 2954 518 2985
rect 552 2954 603 2985
rect 637 2954 688 2988
rect 722 2954 734 2988
rect 334 2948 734 2954
rect -1135 2926 -962 2932
rect -1135 2892 -1123 2926
rect -1089 2892 -1035 2926
rect -1001 2892 -962 2926
rect -1135 2880 -962 2892
rect -910 2880 -877 2932
rect -825 2926 -728 2932
rect -825 2892 -774 2926
rect -740 2892 -728 2926
rect -825 2880 -728 2892
rect -1135 2852 -728 2880
rect -1135 2840 -962 2852
rect -1135 2806 -1123 2840
rect -1089 2806 -1035 2840
rect -1001 2806 -962 2840
rect -1135 2800 -962 2806
rect -910 2800 -877 2852
rect -825 2840 -728 2852
rect -825 2806 -774 2840
rect -740 2806 -728 2840
rect -825 2800 -728 2806
rect 6256 2495 7026 2573
rect 6244 2465 7026 2495
rect 8440 2492 8536 3606
tri 12716 3274 12742 3300 se
rect 12742 3282 13743 3300
tri 13743 3282 13761 3300 sw
rect 12742 3274 13761 3282
rect 12716 3246 13761 3274
rect 12716 3226 12834 3246
tri 12834 3226 12854 3246 nw
tri 13684 3226 13704 3246 ne
rect 10280 3145 10286 3197
rect 10338 3145 10355 3197
rect 10407 3145 10423 3197
rect 10475 3145 10491 3197
rect 10543 3145 10559 3197
rect 10611 3145 10627 3197
rect 10679 3145 10695 3197
rect 10747 3145 10753 3197
rect 12716 3158 12830 3226
tri 12830 3222 12834 3226 nw
rect 10280 3113 10753 3145
rect 10280 3061 10286 3113
rect 10338 3061 10355 3113
rect 10407 3061 10423 3113
rect 10475 3061 10491 3113
rect 10543 3061 10559 3113
rect 10611 3061 10627 3113
rect 10679 3061 10695 3113
rect 10747 3061 10753 3113
rect 13704 2918 13761 3246
tri 13761 2918 13776 2933 sw
rect 9221 2767 9239 2790
rect 12736 2775 12754 2800
rect 16983 2515 17159 3606
rect 23224 3510 23230 3562
rect 23282 3510 23294 3562
rect 23346 3532 24411 3562
tri 24411 3532 24441 3562 sw
rect 23346 3510 24441 3532
tri 24359 3478 24391 3510 ne
rect 22871 3424 22877 3476
rect 22929 3424 22941 3476
rect 22993 3446 24315 3476
tri 24315 3446 24345 3476 sw
rect 22993 3424 24345 3446
tri 24263 3392 24295 3424 ne
rect 24295 3166 24345 3424
rect 24391 3257 24441 3510
tri 24441 3257 24476 3292 sw
rect 24391 3240 24519 3257
tri 24391 3205 24426 3240 ne
rect 24426 3205 24519 3240
rect 24571 3205 24583 3257
rect 24635 3205 24641 3257
tri 24345 3166 24380 3201 sw
rect 24295 3149 24526 3166
tri 24295 3114 24330 3149 ne
rect 24330 3114 24526 3149
rect 24578 3114 24590 3166
rect 24642 3114 24648 3166
rect 24511 3033 24557 3045
rect 24511 2999 24517 3033
rect 24551 2999 24557 3033
rect 24511 2933 24557 2999
rect 24511 2899 24517 2933
rect 24551 2899 24557 2933
rect 23350 2706 23384 2741
rect 24511 2724 24557 2899
rect 24511 2718 24666 2724
rect 24511 2715 24614 2718
rect 24511 2681 24517 2715
rect 24551 2681 24614 2715
rect 24511 2666 24614 2681
rect 24511 2653 24666 2666
rect 24511 2643 24614 2653
rect 24511 2609 24517 2643
rect 24551 2609 24614 2643
rect 24511 2601 24614 2609
rect 24511 2595 24666 2601
rect 15781 2472 15818 2502
rect 6256 2460 7026 2465
rect 18842 2389 19116 2395
rect 18894 2337 18916 2389
rect 18968 2337 18990 2389
rect 19042 2337 19064 2389
rect 18842 2322 19116 2337
rect 18894 2270 18916 2322
rect 18968 2270 18990 2322
rect 19042 2270 19064 2322
rect 18842 2255 19116 2270
rect 18894 2203 18916 2255
rect 18968 2203 18990 2255
rect 19042 2203 19064 2255
rect 18842 2187 19116 2203
rect 18894 2135 18916 2187
rect 18968 2135 18990 2187
rect 19042 2135 19064 2187
rect 18842 2119 19116 2135
rect 18894 2067 18916 2119
rect 18968 2067 18990 2119
rect 19042 2067 19064 2119
rect 18842 2061 19116 2067
rect 20736 2353 20742 2405
rect 20794 2353 20809 2405
rect 20861 2353 20876 2405
rect 20928 2353 20943 2405
rect 20995 2353 21010 2405
rect 21062 2353 21076 2405
rect 21128 2353 21134 2405
rect 20736 2331 21134 2353
rect 20736 2279 20742 2331
rect 20794 2279 20809 2331
rect 20861 2279 20876 2331
rect 20928 2279 20943 2331
rect 20995 2279 21010 2331
rect 21062 2279 21076 2331
rect 21128 2279 21134 2331
rect 22292 2307 22323 2347
rect 20736 2257 21134 2279
rect 20736 2205 20742 2257
rect 20794 2205 20809 2257
rect 20861 2205 20876 2257
rect 20928 2205 20943 2257
rect 20995 2205 21010 2257
rect 21062 2205 21076 2257
rect 21128 2205 21134 2257
rect 20736 2183 21134 2205
rect 20736 2131 20742 2183
rect 20794 2131 20809 2183
rect 20861 2131 20876 2183
rect 20928 2131 20943 2183
rect 20995 2131 21010 2183
rect 21062 2131 21076 2183
rect 21128 2131 21134 2183
rect 20736 2109 21134 2131
rect 20736 2057 20742 2109
rect 20794 2057 20809 2109
rect 20861 2057 20876 2109
rect 20928 2057 20943 2109
rect 20995 2057 21010 2109
rect 21062 2057 21076 2109
rect 21128 2057 21134 2109
rect 10368 1941 10394 1960
rect 12386 1917 12415 1943
rect 10348 1613 10354 1665
rect 10406 1613 10421 1665
rect 10473 1613 10487 1665
rect 10539 1613 10545 1665
rect 10348 1573 10545 1613
rect 10348 1521 10354 1573
rect 10406 1521 10421 1573
rect 10473 1521 10487 1573
rect 10539 1521 10545 1573
rect 24397 1570 24449 1576
rect 24397 1505 24449 1518
rect 24449 1453 24584 1499
rect 24397 1447 24584 1453
rect 24636 1447 24649 1499
rect 24701 1447 24707 1499
rect 25728 1361 25780 1367
tri 25705 1302 25728 1325 se
rect 25728 1302 25780 1309
rect -1144 1299 749 1302
rect -1144 1294 -886 1299
rect -834 1294 -821 1299
rect -769 1294 -756 1299
rect -1144 1260 -1132 1294
rect -1098 1260 -1058 1294
rect -1024 1260 -984 1294
rect -950 1260 -910 1294
rect -769 1260 -762 1294
rect -1144 1247 -886 1260
rect -834 1247 -821 1260
rect -769 1247 -756 1260
rect -704 1247 -691 1299
rect -639 1247 -626 1299
rect -574 1247 -562 1299
rect -510 1294 -498 1299
rect -446 1294 -434 1299
rect -382 1294 -370 1299
rect -318 1294 -306 1299
rect -254 1294 -242 1299
rect -506 1260 -498 1294
rect -254 1260 -246 1294
rect -510 1247 -498 1260
rect -446 1247 -434 1260
rect -382 1247 -370 1260
rect -318 1247 -306 1260
rect -254 1247 -242 1260
rect -190 1247 -178 1299
rect -126 1247 -114 1299
rect -62 1247 -50 1299
rect 2 1294 14 1299
rect 66 1294 78 1299
rect 130 1294 142 1299
rect 194 1294 206 1299
rect 258 1294 270 1299
rect 7 1260 14 1294
rect 258 1260 265 1294
rect 2 1247 14 1260
rect 66 1247 78 1260
rect 130 1247 142 1260
rect 194 1247 206 1260
rect 258 1247 270 1260
rect 322 1247 334 1299
rect 386 1247 398 1299
rect 450 1247 462 1299
rect 514 1294 526 1299
rect 578 1294 590 1299
rect 642 1294 654 1299
rect 706 1294 749 1299
rect 518 1260 526 1294
rect 737 1260 749 1294
tri 25694 1291 25705 1302 se
rect 25705 1297 25780 1302
rect 25705 1291 25728 1297
rect 11939 1264 11976 1289
rect 514 1247 526 1260
rect 578 1247 590 1260
rect 642 1247 654 1260
rect 706 1247 749 1260
rect -1144 1227 749 1247
rect 25095 1239 25101 1291
rect 25153 1239 25165 1291
rect 25217 1245 25728 1291
rect 25217 1239 25780 1245
rect -1144 1220 -886 1227
rect -834 1220 -821 1227
rect -769 1220 -756 1227
rect -1144 1186 -1132 1220
rect -1098 1186 -1058 1220
rect -1024 1186 -984 1220
rect -950 1186 -910 1220
rect -769 1186 -762 1220
rect -1144 1175 -886 1186
rect -834 1175 -821 1186
rect -769 1175 -756 1186
rect -704 1175 -691 1227
rect -639 1175 -626 1227
rect -574 1175 -562 1227
rect -510 1220 -498 1227
rect -446 1220 -434 1227
rect -382 1220 -370 1227
rect -318 1220 -306 1227
rect -254 1220 -242 1227
rect -506 1186 -498 1220
rect -254 1186 -246 1220
rect -510 1175 -498 1186
rect -446 1175 -434 1186
rect -382 1175 -370 1186
rect -318 1175 -306 1186
rect -254 1175 -242 1186
rect -190 1175 -178 1227
rect -126 1175 -114 1227
rect -62 1175 -50 1227
rect 2 1220 14 1227
rect 66 1220 78 1227
rect 130 1220 142 1227
rect 194 1220 206 1227
rect 258 1220 270 1227
rect 7 1186 14 1220
rect 258 1186 265 1220
rect 2 1175 14 1186
rect 66 1175 78 1186
rect 130 1175 142 1186
rect 194 1175 206 1186
rect 258 1175 270 1186
rect 322 1175 334 1227
rect 386 1175 398 1227
rect 450 1175 462 1227
rect 514 1220 526 1227
rect 578 1220 590 1227
rect 642 1220 654 1227
rect 706 1220 749 1227
rect 518 1186 526 1220
rect 737 1186 749 1220
rect 514 1175 526 1186
rect 578 1175 590 1186
rect 642 1175 654 1186
rect 706 1175 749 1186
rect -1144 1155 749 1175
rect -1144 1146 -886 1155
rect -834 1146 -821 1155
rect -769 1146 -756 1155
rect -1144 1112 -1132 1146
rect -1098 1112 -1058 1146
rect -1024 1112 -984 1146
rect -950 1112 -910 1146
rect -769 1112 -762 1146
rect -1144 1103 -886 1112
rect -834 1103 -821 1112
rect -769 1103 -756 1112
rect -704 1103 -691 1155
rect -639 1103 -626 1155
rect -574 1103 -562 1155
rect -510 1146 -498 1155
rect -446 1146 -434 1155
rect -382 1146 -370 1155
rect -318 1146 -306 1155
rect -254 1146 -242 1155
rect -506 1112 -498 1146
rect -254 1112 -246 1146
rect -510 1103 -498 1112
rect -446 1103 -434 1112
rect -382 1103 -370 1112
rect -318 1103 -306 1112
rect -254 1103 -242 1112
rect -190 1103 -178 1155
rect -126 1103 -114 1155
rect -62 1103 -50 1155
rect 2 1146 14 1155
rect 66 1146 78 1155
rect 130 1146 142 1155
rect 194 1146 206 1155
rect 258 1146 270 1155
rect 7 1112 14 1146
rect 258 1112 265 1146
rect 2 1103 14 1112
rect 66 1103 78 1112
rect 130 1103 142 1112
rect 194 1103 206 1112
rect 258 1103 270 1112
rect 322 1103 334 1155
rect 386 1103 398 1155
rect 450 1103 462 1155
rect 514 1146 526 1155
rect 578 1146 590 1155
rect 642 1146 654 1155
rect 706 1146 749 1155
rect 518 1112 526 1146
rect 737 1112 749 1146
rect 23701 1193 25860 1199
rect 23701 1159 23779 1193
rect 23813 1159 23852 1193
rect 23886 1159 23925 1193
rect 23959 1159 23998 1193
rect 24032 1159 24071 1193
rect 24105 1159 24144 1193
rect 24178 1159 24217 1193
rect 24251 1159 24290 1193
rect 24324 1159 24363 1193
rect 24397 1159 24436 1193
rect 24470 1159 24509 1193
rect 24543 1159 24582 1193
rect 24616 1159 24655 1193
rect 24689 1159 24728 1193
rect 24762 1159 24801 1193
rect 24835 1159 24874 1193
rect 24908 1159 24947 1193
rect 24981 1159 25020 1193
rect 25054 1159 25093 1193
rect 25127 1159 25166 1193
rect 25200 1159 25239 1193
rect 25273 1159 25312 1193
rect 25346 1159 25385 1193
rect 25419 1159 25458 1193
rect 25492 1159 25531 1193
rect 25565 1159 25604 1193
rect 25638 1159 25676 1193
rect 25710 1159 25748 1193
rect 25782 1159 25860 1193
rect 23701 1153 25860 1159
rect 514 1103 526 1112
rect 578 1103 590 1112
rect 642 1103 654 1112
rect 706 1103 749 1112
rect -1144 1083 749 1103
rect -1144 1072 -886 1083
rect -834 1072 -821 1083
rect -769 1072 -756 1083
rect -1144 1038 -1132 1072
rect -1098 1038 -1058 1072
rect -1024 1038 -984 1072
rect -950 1038 -910 1072
rect -769 1038 -762 1072
rect -1144 1031 -886 1038
rect -834 1031 -821 1038
rect -769 1031 -756 1038
rect -704 1031 -691 1083
rect -639 1031 -626 1083
rect -574 1031 -562 1083
rect -510 1072 -498 1083
rect -446 1072 -434 1083
rect -382 1072 -370 1083
rect -318 1072 -306 1083
rect -254 1072 -242 1083
rect -506 1038 -498 1072
rect -254 1038 -246 1072
rect -510 1031 -498 1038
rect -446 1031 -434 1038
rect -382 1031 -370 1038
rect -318 1031 -306 1038
rect -254 1031 -242 1038
rect -190 1031 -178 1083
rect -126 1031 -114 1083
rect -62 1031 -50 1083
rect 2 1072 14 1083
rect 66 1072 78 1083
rect 130 1072 142 1083
rect 194 1072 206 1083
rect 258 1072 270 1083
rect 7 1038 14 1072
rect 258 1038 265 1072
rect 2 1031 14 1038
rect 66 1031 78 1038
rect 130 1031 142 1038
rect 194 1031 206 1038
rect 258 1031 270 1038
rect 322 1031 334 1083
rect 386 1031 398 1083
rect 450 1031 462 1083
rect 514 1072 526 1083
rect 578 1072 590 1083
rect 642 1072 654 1083
rect 706 1072 749 1083
rect 518 1038 526 1072
rect 737 1038 749 1072
rect 18784 1126 18964 1132
rect 7822 1038 7857 1068
rect 514 1031 526 1038
rect 578 1031 590 1038
rect 642 1031 654 1038
rect 706 1031 749 1038
rect -1144 1011 749 1031
rect -1144 998 -886 1011
rect -834 998 -821 1011
rect -769 998 -756 1011
rect -1144 964 -1132 998
rect -1098 964 -1058 998
rect -1024 964 -984 998
rect -950 964 -910 998
rect -769 964 -762 998
rect -1144 959 -886 964
rect -834 959 -821 964
rect -769 959 -756 964
rect -704 959 -691 1011
rect -639 959 -626 1011
rect -574 959 -562 1011
rect -510 998 -498 1011
rect -446 998 -434 1011
rect -382 998 -370 1011
rect -318 998 -306 1011
rect -254 998 -242 1011
rect -506 964 -498 998
rect -254 964 -246 998
rect -510 959 -498 964
rect -446 959 -434 964
rect -382 959 -370 964
rect -318 959 -306 964
rect -254 959 -242 964
rect -190 959 -178 1011
rect -126 959 -114 1011
rect -62 959 -50 1011
rect 2 998 14 1011
rect 66 998 78 1011
rect 130 998 142 1011
rect 194 998 206 1011
rect 258 998 270 1011
rect 7 964 14 998
rect 258 964 265 998
rect 2 959 14 964
rect 66 959 78 964
rect 130 959 142 964
rect 194 959 206 964
rect 258 959 270 964
rect 322 959 334 1011
rect 386 959 398 1011
rect 450 959 462 1011
rect 514 998 526 1011
rect 578 998 590 1011
rect 642 998 654 1011
rect 706 998 749 1011
rect 518 964 526 998
rect 737 964 749 998
rect 514 959 526 964
rect 578 959 590 964
rect 642 959 654 964
rect 706 959 749 964
rect -1144 939 749 959
rect 18784 940 18964 946
rect 23701 1121 23749 1153
tri 23749 1121 23781 1153 nw
tri 25780 1121 25812 1153 ne
rect 25812 1121 25860 1153
rect 23701 1120 23748 1121
tri 23748 1120 23749 1121 nw
tri 25812 1120 25813 1121 ne
rect 25813 1120 25820 1121
rect 23701 1105 23747 1120
tri 23747 1119 23748 1120 nw
tri 24748 1119 24749 1120 se
rect 24749 1119 24755 1120
tri 24745 1116 24748 1119 se
rect 24748 1116 24755 1119
rect 23701 1071 23707 1105
rect 23741 1071 23747 1105
rect 23701 979 23747 1071
rect 24414 1110 24755 1116
rect 24414 1076 24426 1110
rect 24460 1076 24500 1110
rect 24534 1076 24574 1110
rect 24608 1076 24648 1110
rect 24682 1076 24755 1110
rect 24414 1070 24755 1076
tri 24747 1068 24749 1070 ne
rect 24749 1068 24755 1070
rect 24807 1068 24819 1120
rect 24871 1119 24877 1120
tri 24877 1119 24878 1120 sw
tri 25813 1119 25814 1120 ne
rect 24871 1116 24878 1119
tri 24878 1116 24881 1119 sw
rect 24871 1110 25454 1116
rect 24871 1076 25186 1110
rect 25220 1076 25260 1110
rect 25294 1076 25334 1110
rect 25368 1076 25408 1110
rect 25442 1076 25454 1110
rect 24871 1070 25454 1076
rect 25814 1087 25820 1120
rect 25854 1087 25860 1121
rect 24871 1068 24877 1070
tri 24877 1068 24879 1070 nw
rect 25814 1042 25860 1087
rect 23948 989 23954 1041
rect 24006 989 24019 1041
rect 24071 1035 24077 1041
tri 24077 1035 24083 1041 sw
rect 24071 1029 25130 1035
rect 24071 995 24130 1029
rect 24164 995 24229 1029
rect 24263 995 24328 1029
rect 24362 995 24899 1029
rect 24933 995 24992 1029
rect 25026 995 25084 1029
rect 25118 995 25130 1029
rect 24071 989 25130 995
rect 25814 1008 25820 1042
rect 25854 1008 25860 1042
rect 23701 945 23707 979
rect 23741 945 23747 979
tri 25551 972 25563 984 se
rect 25563 972 25609 984
tri 25540 961 25551 972 se
rect 25551 961 25569 972
rect -1144 924 -886 939
rect -834 924 -821 939
rect -769 924 -756 939
rect -1144 890 -1132 924
rect -1098 890 -1058 924
rect -1024 890 -984 924
rect -950 890 -910 924
rect -769 890 -762 924
rect -1144 887 -886 890
rect -834 887 -821 890
rect -769 887 -756 890
rect -704 887 -691 939
rect -639 887 -626 939
rect -574 887 -562 939
rect -510 924 -498 939
rect -446 924 -434 939
rect -382 924 -370 939
rect -318 924 -306 939
rect -254 924 -242 939
rect -506 890 -498 924
rect -254 890 -246 924
rect -510 887 -498 890
rect -446 887 -434 890
rect -382 887 -370 890
rect -318 887 -306 890
rect -254 887 -242 890
rect -190 887 -178 939
rect -126 887 -114 939
rect -62 887 -50 939
rect 2 924 14 939
rect 66 924 78 939
rect 130 924 142 939
rect 194 924 206 939
rect 258 924 270 939
rect 7 890 14 924
rect 258 890 265 924
rect 2 887 14 890
rect 66 887 78 890
rect 130 887 142 890
rect 194 887 206 890
rect 258 887 270 890
rect 322 887 334 939
rect 386 887 398 939
rect 450 887 462 939
rect 514 924 526 939
rect 578 924 590 939
rect 642 924 654 939
rect 706 924 749 939
rect 518 890 526 924
rect 737 890 749 924
rect 514 887 526 890
rect 578 887 590 890
rect 642 887 654 890
rect 706 887 749 890
rect -1144 867 749 887
rect -1144 850 -886 867
rect -834 850 -821 867
rect -769 850 -756 867
rect -1144 816 -1132 850
rect -1098 816 -1058 850
rect -1024 816 -984 850
rect -950 816 -910 850
rect -769 816 -762 850
rect -1144 815 -886 816
rect -834 815 -821 816
rect -769 815 -756 816
rect -704 815 -691 867
rect -639 815 -626 867
rect -574 815 -562 867
rect -510 850 -498 867
rect -446 850 -434 867
rect -382 850 -370 867
rect -318 850 -306 867
rect -254 850 -242 867
rect -506 816 -498 850
rect -254 816 -246 850
rect -510 815 -498 816
rect -446 815 -434 816
rect -382 815 -370 816
rect -318 815 -306 816
rect -254 815 -242 816
rect -190 815 -178 867
rect -126 815 -114 867
rect -62 815 -50 867
rect 2 850 14 867
rect 66 850 78 867
rect 130 850 142 867
rect 194 850 206 867
rect 258 850 270 867
rect 7 816 14 850
rect 258 816 265 850
rect 2 815 14 816
rect 66 815 78 816
rect 130 815 142 816
rect 194 815 206 816
rect 258 815 270 816
rect 322 815 334 867
rect 386 815 398 867
rect 450 815 462 867
rect 514 850 526 867
rect 578 850 590 867
rect 642 850 654 867
rect 706 850 749 867
rect 518 816 526 850
rect 737 816 749 850
rect 514 815 526 816
rect 578 815 590 816
rect 642 815 654 816
rect 706 815 749 816
rect -1144 808 749 815
rect 23701 893 23747 945
rect 23701 859 23707 893
rect 23741 859 23747 893
rect -1144 807 712 808
rect 23701 807 23747 859
rect 23947 945 23993 957
rect 23947 911 23953 945
rect 23987 911 23993 945
tri 24048 940 24051 943 se
rect 24051 940 24057 943
rect 23947 873 23993 911
rect 24044 934 24057 940
rect 24044 900 24056 934
rect 24044 894 24057 900
tri 24048 891 24051 894 ne
rect 24051 891 24057 894
rect 24109 891 24121 943
rect 24173 891 24179 943
tri 24335 940 24337 942 se
rect 24337 940 24343 943
rect 24335 894 24343 940
tri 24335 892 24337 894 ne
rect 24337 891 24343 894
rect 24395 891 24407 943
rect 24459 891 24465 943
rect 24618 891 24624 943
rect 24676 891 24688 943
rect 24740 940 24746 943
tri 24746 940 24748 942 sw
rect 24740 894 24748 940
rect 24740 891 24746 894
tri 24746 892 24748 894 nw
rect 24823 906 24869 918
rect 23947 839 23953 873
rect 23987 872 23993 873
tri 23993 872 23997 876 sw
rect 24823 872 24829 906
rect 24863 872 24869 906
rect 24925 909 24931 961
rect 24983 909 24995 961
rect 25047 938 25569 961
rect 25603 938 25609 972
rect 25047 933 25609 938
rect 25047 929 25085 933
tri 25085 929 25089 933 nw
tri 25231 929 25235 933 ne
rect 25235 929 25425 933
tri 25425 929 25429 933 nw
tri 25529 929 25533 933 ne
rect 25533 929 25609 933
rect 25047 927 25083 929
tri 25083 927 25085 929 nw
tri 25235 927 25237 929 ne
rect 25237 927 25413 929
rect 25047 909 25055 927
rect 24925 893 24937 909
rect 24971 893 25009 909
rect 25043 893 25055 909
tri 25055 899 25083 927 nw
tri 25237 899 25265 927 ne
rect 24925 887 25055 893
rect 23987 859 23997 872
tri 23997 859 24010 872 sw
rect 23987 856 24010 859
tri 24010 856 24013 859 sw
rect 23987 850 24013 856
tri 24013 850 24019 856 sw
rect 23987 842 24019 850
tri 24019 842 24027 850 sw
rect 24823 847 24869 872
tri 24869 847 24872 850 sw
rect 25095 847 25101 899
rect 25153 847 25165 899
rect 25217 853 25225 899
rect 25265 893 25277 927
rect 25311 893 25349 927
rect 25383 917 25413 927
tri 25413 917 25425 929 nw
tri 25533 917 25545 929 ne
rect 25545 917 25609 929
rect 25814 963 25860 1008
rect 25814 929 25820 963
rect 25854 929 25860 963
rect 25383 902 25398 917
tri 25398 902 25413 917 nw
tri 25545 902 25560 917 ne
rect 25560 902 25609 917
rect 25383 900 25396 902
tri 25396 900 25398 902 nw
rect 25383 893 25395 900
tri 25395 899 25396 900 nw
rect 25265 887 25395 893
rect 25447 890 25493 902
tri 25560 900 25562 902 ne
rect 25562 900 25609 902
tri 25562 899 25563 900 ne
rect 25217 847 25223 853
tri 25223 851 25225 853 nw
rect 25447 856 25453 890
rect 25487 856 25493 890
tri 25444 847 25447 850 se
rect 25447 847 25493 856
rect 25563 866 25569 900
rect 25603 866 25609 900
rect 25563 854 25609 866
rect 25645 911 25697 917
rect 23987 839 24780 842
rect 23947 836 24780 839
rect 23947 814 24215 836
tri 23382 773 23397 788 se
tri 23380 771 23382 773 se
rect 23382 771 23397 773
tri 23363 754 23380 771 se
rect 23380 754 23397 771
rect 23701 773 23707 807
rect 23741 773 23747 807
tri 24185 802 24197 814 ne
rect 24197 802 24215 814
rect 24249 802 24287 836
rect 24321 814 24477 836
rect 24321 802 24339 814
tri 24339 802 24351 814 nw
tri 24447 802 24459 814 ne
rect 24459 802 24477 814
rect 24511 802 24549 836
rect 24583 814 24780 836
rect 24583 802 24599 814
tri 24197 800 24199 802 ne
rect 24199 800 24337 802
tri 24337 800 24339 802 nw
tri 24459 800 24461 802 ne
rect 24461 800 24599 802
tri 24599 800 24613 814 nw
tri 24700 800 24714 814 ne
rect 24714 800 24780 814
tri 24199 796 24203 800 ne
rect 24203 796 24333 800
tri 24333 796 24337 800 nw
tri 24461 796 24465 800 ne
rect 24465 796 24595 800
tri 24595 796 24599 800 nw
tri 24714 796 24718 800 ne
rect 24718 796 24780 800
tri 24718 784 24730 796 ne
rect 24730 784 24780 796
rect 24823 834 24872 847
rect 24823 800 24829 834
rect 24863 818 24872 834
tri 24872 818 24901 847 sw
tri 25415 818 25444 847 se
rect 25444 818 25493 847
rect 24863 816 24901 818
tri 24901 816 24903 818 sw
tri 25413 816 25415 818 se
rect 25415 816 25453 818
rect 24863 800 25453 816
rect 24823 788 25453 800
tri 25431 784 25435 788 ne
rect 25435 784 25453 788
rect 25487 816 25493 818
tri 25493 816 25527 850 sw
tri 25611 816 25645 850 se
rect 25645 847 25697 859
rect 25487 795 25645 816
rect 25487 789 25697 795
rect 25814 884 25860 929
rect 25814 850 25820 884
rect 25854 850 25860 884
rect 25814 805 25860 850
rect 25487 788 25695 789
rect 25487 784 25493 788
tri 24730 780 24734 784 ne
rect 23701 721 23747 773
rect 24734 741 24780 784
tri 25435 772 25447 784 ne
rect 25447 772 25493 784
tri 25493 772 25509 788 nw
rect 25814 771 25820 805
rect 25854 771 25860 805
tri 24780 741 24799 760 sw
rect 24734 740 24833 741
tri 24734 727 24747 740 ne
rect 24747 727 24833 740
tri 23384 703 23397 716 ne
rect 23701 687 23707 721
rect 23741 687 23747 721
tri 24747 693 24781 727 ne
rect 24781 693 24833 727
tri 24781 689 24785 693 ne
rect 24785 689 24833 693
rect 24885 689 24897 741
rect 24949 689 24955 741
rect 25814 727 25860 771
rect 25814 693 25820 727
rect 25854 693 25860 727
rect 23701 655 23747 687
tri 23747 655 23781 689 sw
tri 25780 655 25814 689 se
rect 25814 655 25860 693
rect 23701 649 25860 655
tri 23034 615 23064 645 ne
rect 23064 615 23068 645
tri 23064 611 23068 615 ne
rect 23701 615 23779 649
rect 23813 615 23851 649
rect 23885 615 23923 649
rect 23957 615 23996 649
rect 24030 615 24069 649
rect 24103 615 24142 649
rect 24176 615 24215 649
rect 24249 615 24288 649
rect 24322 615 24361 649
rect 24395 615 24434 649
rect 24468 615 24501 649
rect 24553 615 24580 649
rect 24614 615 24653 649
rect 24687 615 24726 649
rect 24760 615 24799 649
rect 24833 615 24872 649
rect 24906 615 24945 649
rect 24979 615 25018 649
rect 25052 615 25091 649
rect 25125 615 25164 649
rect 25198 615 25237 649
rect 25271 615 25310 649
rect 25344 615 25383 649
rect 25417 615 25456 649
rect 25490 615 25529 649
rect 25563 615 25602 649
rect 25636 615 25675 649
rect 25709 615 25748 649
rect 25782 615 25860 649
rect 23701 609 24501 615
tri 24467 575 24501 609 ne
rect 24553 609 25860 615
rect 24501 563 24553 597
tri 24553 575 24587 609 nw
tri 23253 522 23277 546 se
rect 23277 522 23283 546
tri 22873 509 22886 522 se
rect 22886 509 23283 522
tri 12307 494 12322 509 sw
tri 22858 494 22873 509 se
rect 22873 494 23283 509
rect 23335 494 23347 546
rect 23399 494 23405 546
rect 24501 505 24553 511
rect 12307 438 12322 494
tri 12322 438 12378 494 sw
tri 22839 475 22858 494 se
rect 22858 475 22881 494
tri 22881 475 22900 494 nw
tri 22802 438 22839 475 se
rect 22839 438 22844 475
tri 22844 438 22881 475 nw
tri 23028 440 23031 443 sw
rect 12307 321 13506 438
tri 22797 433 22802 438 se
rect 22802 433 22839 438
tri 22839 433 22844 438 nw
tri 22783 419 22797 433 se
rect 22797 419 22825 433
tri 22825 419 22839 433 nw
rect 22418 391 22797 419
tri 22797 391 22825 419 nw
tri 23028 397 23031 400 nw
rect 22418 346 22446 391
tri 22986 361 22992 367 se
tri 13124 281 13164 321 ne
rect 13164 281 13506 321
tri 20449 318 20477 346 se
rect 20477 318 22446 346
tri 20448 317 20449 318 se
rect 20449 317 20489 318
tri 20489 317 20490 318 nw
tri 20412 281 20448 317 se
rect 20448 281 20453 317
tri 20453 281 20489 317 nw
tri 13164 229 13216 281 ne
rect 13216 258 13506 281
tri 13506 258 13529 281 sw
tri 20407 276 20412 281 se
rect 20412 276 20448 281
tri 20448 276 20453 281 nw
tri 20389 258 20407 276 se
rect 20407 258 20430 276
tri 20430 258 20448 276 nw
rect 13216 229 13529 258
tri 13529 229 13558 258 sw
tri 16091 229 16120 258 se
rect 16120 229 16412 258
tri 20366 235 20389 258 se
rect 20389 235 20407 258
tri 20407 235 20430 258 nw
rect -253 225 -247 229
rect -730 219 -247 225
rect -678 197 -247 219
rect -253 177 -247 197
rect -195 177 -183 229
rect -131 177 -125 229
tri 13216 214 13231 229 ne
rect 13231 208 13558 229
tri 13558 208 13579 229 sw
tri 16070 208 16091 229 se
rect 16091 208 16412 229
rect -730 155 -678 167
rect -730 97 -678 103
rect 13231 154 16412 208
tri 20325 194 20366 235 se
tri 20366 194 20407 235 nw
tri 20312 181 20325 194 se
rect 20325 181 20353 194
tri 20353 181 20366 194 nw
rect 13231 129 13852 154
tri 13852 129 13877 154 nw
rect 19407 129 19413 181
rect 19465 129 19477 181
rect 19529 153 20325 181
tri 20325 153 20353 181 nw
rect 19529 129 19535 153
rect 13231 -13 13829 129
tri 13829 106 13852 129 nw
rect 13231 -65 13237 -13
rect 13289 -65 13304 -13
rect 13356 -65 13371 -13
rect 13423 -65 13438 -13
rect 13490 -65 13505 -13
rect 13557 -65 13572 -13
rect 13624 -65 13639 -13
rect 13691 -65 13705 -13
rect 13757 -65 13771 -13
rect 13823 -65 13829 -13
rect 13231 -117 13829 -65
rect 13231 -169 13237 -117
rect 13289 -169 13304 -117
rect 13356 -169 13371 -117
rect 13423 -169 13438 -117
rect 13490 -169 13505 -117
rect 13557 -169 13572 -117
rect 13624 -169 13639 -117
rect 13691 -169 13705 -117
rect 13757 -169 13771 -117
rect 13823 -169 13829 -117
rect -613 -3123 -582 -3083
rect -369 -4361 766 -4345
rect -369 -4413 641 -4361
rect 693 -4413 707 -4361
rect 759 -4413 766 -4361
rect -369 -4430 766 -4413
rect -286 -4433 -251 -4430
rect -803 -5553 -780 -5527
rect -1112 -6297 -1047 -6246
rect 707 -6388 744 -6358
rect -294 -6430 -277 -6408
<< via1 >>
rect 1357 22393 1409 22407
rect 1357 22359 1366 22393
rect 1366 22359 1400 22393
rect 1400 22359 1409 22393
rect 1357 22355 1409 22359
rect 1357 22321 1409 22343
rect 1357 22291 1366 22321
rect 1366 22291 1400 22321
rect 1400 22291 1409 22321
rect 1513 22393 1565 22407
rect 1513 22359 1522 22393
rect 1522 22359 1556 22393
rect 1556 22359 1565 22393
rect 1513 22355 1565 22359
rect 1513 22321 1565 22343
rect 1513 22291 1522 22321
rect 1522 22291 1556 22321
rect 1556 22291 1565 22321
rect 1435 22221 1444 22245
rect 1444 22221 1478 22245
rect 1478 22221 1487 22245
rect 1435 22193 1487 22221
rect 1435 22149 1444 22181
rect 1444 22149 1478 22181
rect 1478 22149 1487 22181
rect 1435 22129 1487 22149
rect 1435 22111 1487 22117
rect 1435 22077 1444 22111
rect 1444 22077 1478 22111
rect 1478 22077 1487 22111
rect 1435 22065 1487 22077
rect 1279 21895 1331 21907
rect 1279 21861 1288 21895
rect 1288 21861 1322 21895
rect 1322 21861 1331 21895
rect 1279 21855 1331 21861
rect 1279 21823 1331 21843
rect 1279 21791 1288 21823
rect 1288 21791 1322 21823
rect 1322 21791 1331 21823
rect 1279 21751 1331 21779
rect 1279 21727 1288 21751
rect 1288 21727 1322 21751
rect 1322 21727 1331 21751
rect 1591 21895 1643 21907
rect 1591 21861 1600 21895
rect 1600 21861 1634 21895
rect 1634 21861 1643 21895
rect 1591 21855 1643 21861
rect 1591 21823 1643 21843
rect 1591 21791 1600 21823
rect 1600 21791 1634 21823
rect 1634 21791 1643 21823
rect 1591 21751 1643 21779
rect 1591 21727 1600 21751
rect 1600 21727 1634 21751
rect 1634 21727 1643 21751
rect 1279 21559 1288 21583
rect 1288 21559 1322 21583
rect 1322 21559 1331 21583
rect 1279 21531 1331 21559
rect 1279 21487 1288 21519
rect 1288 21487 1322 21519
rect 1322 21487 1331 21519
rect 1279 21467 1331 21487
rect 1279 21449 1331 21455
rect 1279 21415 1288 21449
rect 1288 21415 1322 21449
rect 1322 21415 1331 21449
rect 1279 21403 1331 21415
rect 1591 21559 1600 21583
rect 1600 21559 1634 21583
rect 1634 21559 1643 21583
rect 1591 21531 1643 21559
rect 1591 21487 1600 21519
rect 1600 21487 1634 21519
rect 1634 21487 1643 21519
rect 1591 21467 1643 21487
rect 1591 21449 1643 21455
rect 1591 21415 1600 21449
rect 1600 21415 1634 21449
rect 1634 21415 1643 21449
rect 1591 21403 1643 21415
rect 1435 21233 1487 21245
rect 1435 21199 1444 21233
rect 1444 21199 1478 21233
rect 1478 21199 1487 21233
rect 1435 21193 1487 21199
rect 1435 21161 1487 21181
rect 1435 21129 1444 21161
rect 1444 21129 1478 21161
rect 1478 21129 1487 21161
rect 1435 21089 1487 21117
rect 1435 21065 1444 21089
rect 1444 21065 1478 21089
rect 1478 21065 1487 21089
rect 2020 14588 2072 14640
rect 2020 14513 2072 14565
rect 2112 14588 2164 14640
rect 2112 14513 2164 14565
rect 1341 14250 1393 14302
rect 1341 14175 1393 14227
rect 1433 14248 1485 14300
rect 1433 14173 1485 14225
rect 1341 10704 1393 10756
rect 1678 10704 1730 10756
rect 1341 10637 1393 10689
rect 1678 10637 1730 10689
rect 1678 10499 1730 10505
rect 1678 10465 1687 10499
rect 1687 10465 1721 10499
rect 1721 10465 1730 10499
rect 1678 10453 1730 10465
rect 1678 10426 1730 10435
rect 1678 10392 1687 10426
rect 1687 10392 1721 10426
rect 1721 10392 1730 10426
rect 2419 10489 2471 10541
rect 2419 10425 2471 10477
rect 1678 10383 1730 10392
rect 1678 10352 1730 10364
rect 1678 10318 1687 10352
rect 1687 10318 1721 10352
rect 1721 10318 1730 10352
rect 1678 10312 1730 10318
rect 1163 10022 1215 10074
rect 1163 9958 1215 10010
rect 2171 10022 2223 10074
rect 2171 9958 2223 10010
rect 2419 9818 2471 9870
rect 2419 9754 2471 9806
rect 1433 9645 1485 9697
rect 1433 9575 1485 9627
rect 1433 9504 1485 9556
rect 2337 9462 2389 9514
rect 1163 9408 1215 9460
rect 1163 9344 1215 9396
rect 2337 9398 2389 9450
rect 25526 6336 25578 6388
rect 25590 6336 25642 6388
rect 2100 6281 2152 6333
rect 2164 6281 2216 6333
rect 1932 6207 1984 6259
rect 1996 6207 2048 6259
rect 25069 6241 25121 6293
rect 25133 6241 25185 6293
rect 2255 5936 2307 5988
rect 2255 5872 2307 5924
rect 8667 5941 8719 5993
rect 8731 5941 8783 5993
rect 2359 5866 2411 5918
rect 2423 5866 2475 5918
rect 13064 5866 13116 5918
rect 13128 5866 13180 5918
rect 7348 5149 7400 5201
rect 7412 5149 7464 5201
rect 7888 5149 7940 5201
rect 7952 5149 8004 5201
rect 25416 5184 25468 5236
rect 25325 5124 25377 5176
rect 25416 5104 25468 5156
rect 25325 5044 25377 5096
rect -962 3040 -910 3092
rect -877 3040 -825 3092
rect -962 2960 -910 3012
rect -877 2960 -825 3012
rect -617 3032 -585 3056
rect -585 3032 -565 3056
rect -617 3004 -565 3032
rect -535 3032 -533 3056
rect -533 3032 -499 3056
rect -499 3032 -483 3056
rect -535 3004 -483 3032
rect -453 3032 -447 3056
rect -447 3032 -413 3056
rect -413 3032 -401 3056
rect -453 3004 -401 3032
rect -371 3032 -362 3056
rect -362 3032 -328 3056
rect -328 3032 -319 3056
rect -371 3004 -319 3032
rect -289 3032 -277 3056
rect -277 3032 -243 3056
rect -243 3032 -237 3056
rect -289 3004 -237 3032
rect -141 3032 -139 3037
rect -139 3032 -105 3037
rect -105 3032 -89 3037
rect -141 2988 -89 3032
rect -141 2985 -139 2988
rect -139 2985 -105 2988
rect -105 2985 -89 2988
rect -65 3032 -53 3037
rect -53 3032 -19 3037
rect -19 3032 -13 3037
rect -65 2988 -13 3032
rect -65 2985 -53 2988
rect -53 2985 -19 2988
rect -19 2985 -13 2988
rect 11 3032 33 3037
rect 33 3032 63 3037
rect 86 3032 118 3037
rect 118 3032 138 3037
rect 11 2988 63 3032
rect 86 2988 138 3032
rect 11 2985 33 2988
rect 33 2985 63 2988
rect 86 2985 118 2988
rect 118 2985 138 2988
rect 357 3032 380 3037
rect 380 3032 409 3037
rect 433 3032 466 3037
rect 466 3032 485 3037
rect 357 2988 409 3032
rect 433 2988 485 3032
rect 357 2985 380 2988
rect 380 2985 409 2988
rect 433 2985 466 2988
rect 466 2985 485 2988
rect 509 3032 518 3037
rect 518 3032 552 3037
rect 552 3032 561 3037
rect 509 2988 561 3032
rect 509 2985 518 2988
rect 518 2985 552 2988
rect 552 2985 561 2988
rect 584 3032 603 3037
rect 603 3032 636 3037
rect 584 2988 636 3032
rect 584 2985 603 2988
rect 603 2985 636 2988
rect -962 2926 -910 2932
rect -962 2892 -948 2926
rect -948 2892 -914 2926
rect -914 2892 -910 2926
rect -962 2880 -910 2892
rect -877 2926 -825 2932
rect -877 2892 -861 2926
rect -861 2892 -827 2926
rect -827 2892 -825 2926
rect -877 2880 -825 2892
rect -962 2840 -910 2852
rect -962 2806 -948 2840
rect -948 2806 -914 2840
rect -914 2806 -910 2840
rect -962 2800 -910 2806
rect -877 2840 -825 2852
rect -877 2806 -861 2840
rect -861 2806 -827 2840
rect -827 2806 -825 2840
rect -877 2800 -825 2806
rect 10286 3145 10338 3197
rect 10355 3145 10407 3197
rect 10423 3145 10475 3197
rect 10491 3145 10543 3197
rect 10559 3145 10611 3197
rect 10627 3145 10679 3197
rect 10695 3145 10747 3197
rect 10286 3061 10338 3113
rect 10355 3061 10407 3113
rect 10423 3061 10475 3113
rect 10491 3061 10543 3113
rect 10559 3061 10611 3113
rect 10627 3061 10679 3113
rect 10695 3061 10747 3113
rect 23230 3510 23282 3562
rect 23294 3510 23346 3562
rect 22877 3424 22929 3476
rect 22941 3424 22993 3476
rect 24519 3205 24571 3257
rect 24583 3205 24635 3257
rect 24526 3114 24578 3166
rect 24590 3114 24642 3166
rect 24614 2666 24666 2718
rect 24614 2601 24666 2653
rect 18842 2337 18894 2389
rect 18916 2337 18968 2389
rect 18990 2337 19042 2389
rect 19064 2337 19116 2389
rect 18842 2270 18894 2322
rect 18916 2270 18968 2322
rect 18990 2270 19042 2322
rect 19064 2270 19116 2322
rect 18842 2203 18894 2255
rect 18916 2203 18968 2255
rect 18990 2203 19042 2255
rect 19064 2203 19116 2255
rect 18842 2135 18894 2187
rect 18916 2135 18968 2187
rect 18990 2135 19042 2187
rect 19064 2135 19116 2187
rect 18842 2067 18894 2119
rect 18916 2067 18968 2119
rect 18990 2067 19042 2119
rect 19064 2067 19116 2119
rect 20742 2353 20794 2405
rect 20809 2353 20861 2405
rect 20876 2353 20928 2405
rect 20943 2353 20995 2405
rect 21010 2353 21062 2405
rect 21076 2353 21128 2405
rect 20742 2279 20794 2331
rect 20809 2279 20861 2331
rect 20876 2279 20928 2331
rect 20943 2279 20995 2331
rect 21010 2279 21062 2331
rect 21076 2279 21128 2331
rect 20742 2205 20794 2257
rect 20809 2205 20861 2257
rect 20876 2205 20928 2257
rect 20943 2205 20995 2257
rect 21010 2205 21062 2257
rect 21076 2205 21128 2257
rect 20742 2131 20794 2183
rect 20809 2131 20861 2183
rect 20876 2131 20928 2183
rect 20943 2131 20995 2183
rect 21010 2131 21062 2183
rect 21076 2131 21128 2183
rect 20742 2057 20794 2109
rect 20809 2057 20861 2109
rect 20876 2057 20928 2109
rect 20943 2057 20995 2109
rect 21010 2057 21062 2109
rect 21076 2057 21128 2109
rect 10354 1613 10406 1665
rect 10421 1613 10473 1665
rect 10487 1613 10539 1665
rect 10354 1521 10406 1573
rect 10421 1521 10473 1573
rect 10487 1521 10539 1573
rect 24397 1518 24449 1570
rect 24397 1453 24449 1505
rect 24584 1447 24636 1499
rect 24649 1447 24701 1499
rect 25728 1309 25780 1361
rect -886 1294 -834 1299
rect -821 1294 -769 1299
rect -756 1294 -704 1299
rect -886 1260 -876 1294
rect -876 1260 -836 1294
rect -836 1260 -834 1294
rect -821 1260 -802 1294
rect -802 1260 -769 1294
rect -756 1260 -728 1294
rect -728 1260 -704 1294
rect -886 1247 -834 1260
rect -821 1247 -769 1260
rect -756 1247 -704 1260
rect -691 1294 -639 1299
rect -691 1260 -688 1294
rect -688 1260 -654 1294
rect -654 1260 -639 1294
rect -691 1247 -639 1260
rect -626 1294 -574 1299
rect -626 1260 -614 1294
rect -614 1260 -580 1294
rect -580 1260 -574 1294
rect -626 1247 -574 1260
rect -562 1294 -510 1299
rect -498 1294 -446 1299
rect -434 1294 -382 1299
rect -370 1294 -318 1299
rect -306 1294 -254 1299
rect -242 1294 -190 1299
rect -562 1260 -540 1294
rect -540 1260 -510 1294
rect -498 1260 -466 1294
rect -466 1260 -446 1294
rect -434 1260 -432 1294
rect -432 1260 -392 1294
rect -392 1260 -382 1294
rect -370 1260 -358 1294
rect -358 1260 -319 1294
rect -319 1260 -318 1294
rect -306 1260 -285 1294
rect -285 1260 -254 1294
rect -242 1260 -212 1294
rect -212 1260 -190 1294
rect -562 1247 -510 1260
rect -498 1247 -446 1260
rect -434 1247 -382 1260
rect -370 1247 -318 1260
rect -306 1247 -254 1260
rect -242 1247 -190 1260
rect -178 1294 -126 1299
rect -178 1260 -173 1294
rect -173 1260 -139 1294
rect -139 1260 -126 1294
rect -178 1247 -126 1260
rect -114 1294 -62 1299
rect -114 1260 -100 1294
rect -100 1260 -66 1294
rect -66 1260 -62 1294
rect -114 1247 -62 1260
rect -50 1294 2 1299
rect 14 1294 66 1299
rect 78 1294 130 1299
rect 142 1294 194 1299
rect 206 1294 258 1299
rect 270 1294 322 1299
rect -50 1260 -27 1294
rect -27 1260 2 1294
rect 14 1260 46 1294
rect 46 1260 66 1294
rect 78 1260 80 1294
rect 80 1260 119 1294
rect 119 1260 130 1294
rect 142 1260 153 1294
rect 153 1260 192 1294
rect 192 1260 194 1294
rect 206 1260 226 1294
rect 226 1260 258 1294
rect 270 1260 299 1294
rect 299 1260 322 1294
rect -50 1247 2 1260
rect 14 1247 66 1260
rect 78 1247 130 1260
rect 142 1247 194 1260
rect 206 1247 258 1260
rect 270 1247 322 1260
rect 334 1294 386 1299
rect 334 1260 338 1294
rect 338 1260 372 1294
rect 372 1260 386 1294
rect 334 1247 386 1260
rect 398 1294 450 1299
rect 398 1260 411 1294
rect 411 1260 445 1294
rect 445 1260 450 1294
rect 398 1247 450 1260
rect 462 1294 514 1299
rect 526 1294 578 1299
rect 590 1294 642 1299
rect 654 1294 706 1299
rect 462 1260 484 1294
rect 484 1260 514 1294
rect 526 1260 557 1294
rect 557 1260 578 1294
rect 590 1260 591 1294
rect 591 1260 630 1294
rect 630 1260 642 1294
rect 654 1260 664 1294
rect 664 1260 703 1294
rect 703 1260 706 1294
rect 462 1247 514 1260
rect 526 1247 578 1260
rect 590 1247 642 1260
rect 654 1247 706 1260
rect 25101 1239 25153 1291
rect 25165 1239 25217 1291
rect 25728 1245 25780 1297
rect -886 1220 -834 1227
rect -821 1220 -769 1227
rect -756 1220 -704 1227
rect -886 1186 -876 1220
rect -876 1186 -836 1220
rect -836 1186 -834 1220
rect -821 1186 -802 1220
rect -802 1186 -769 1220
rect -756 1186 -728 1220
rect -728 1186 -704 1220
rect -886 1175 -834 1186
rect -821 1175 -769 1186
rect -756 1175 -704 1186
rect -691 1220 -639 1227
rect -691 1186 -688 1220
rect -688 1186 -654 1220
rect -654 1186 -639 1220
rect -691 1175 -639 1186
rect -626 1220 -574 1227
rect -626 1186 -614 1220
rect -614 1186 -580 1220
rect -580 1186 -574 1220
rect -626 1175 -574 1186
rect -562 1220 -510 1227
rect -498 1220 -446 1227
rect -434 1220 -382 1227
rect -370 1220 -318 1227
rect -306 1220 -254 1227
rect -242 1220 -190 1227
rect -562 1186 -540 1220
rect -540 1186 -510 1220
rect -498 1186 -466 1220
rect -466 1186 -446 1220
rect -434 1186 -432 1220
rect -432 1186 -392 1220
rect -392 1186 -382 1220
rect -370 1186 -358 1220
rect -358 1186 -319 1220
rect -319 1186 -318 1220
rect -306 1186 -285 1220
rect -285 1186 -254 1220
rect -242 1186 -212 1220
rect -212 1186 -190 1220
rect -562 1175 -510 1186
rect -498 1175 -446 1186
rect -434 1175 -382 1186
rect -370 1175 -318 1186
rect -306 1175 -254 1186
rect -242 1175 -190 1186
rect -178 1220 -126 1227
rect -178 1186 -173 1220
rect -173 1186 -139 1220
rect -139 1186 -126 1220
rect -178 1175 -126 1186
rect -114 1220 -62 1227
rect -114 1186 -100 1220
rect -100 1186 -66 1220
rect -66 1186 -62 1220
rect -114 1175 -62 1186
rect -50 1220 2 1227
rect 14 1220 66 1227
rect 78 1220 130 1227
rect 142 1220 194 1227
rect 206 1220 258 1227
rect 270 1220 322 1227
rect -50 1186 -27 1220
rect -27 1186 2 1220
rect 14 1186 46 1220
rect 46 1186 66 1220
rect 78 1186 80 1220
rect 80 1186 119 1220
rect 119 1186 130 1220
rect 142 1186 153 1220
rect 153 1186 192 1220
rect 192 1186 194 1220
rect 206 1186 226 1220
rect 226 1186 258 1220
rect 270 1186 299 1220
rect 299 1186 322 1220
rect -50 1175 2 1186
rect 14 1175 66 1186
rect 78 1175 130 1186
rect 142 1175 194 1186
rect 206 1175 258 1186
rect 270 1175 322 1186
rect 334 1220 386 1227
rect 334 1186 338 1220
rect 338 1186 372 1220
rect 372 1186 386 1220
rect 334 1175 386 1186
rect 398 1220 450 1227
rect 398 1186 411 1220
rect 411 1186 445 1220
rect 445 1186 450 1220
rect 398 1175 450 1186
rect 462 1220 514 1227
rect 526 1220 578 1227
rect 590 1220 642 1227
rect 654 1220 706 1227
rect 462 1186 484 1220
rect 484 1186 514 1220
rect 526 1186 557 1220
rect 557 1186 578 1220
rect 590 1186 591 1220
rect 591 1186 630 1220
rect 630 1186 642 1220
rect 654 1186 664 1220
rect 664 1186 703 1220
rect 703 1186 706 1220
rect 462 1175 514 1186
rect 526 1175 578 1186
rect 590 1175 642 1186
rect 654 1175 706 1186
rect -886 1146 -834 1155
rect -821 1146 -769 1155
rect -756 1146 -704 1155
rect -886 1112 -876 1146
rect -876 1112 -836 1146
rect -836 1112 -834 1146
rect -821 1112 -802 1146
rect -802 1112 -769 1146
rect -756 1112 -728 1146
rect -728 1112 -704 1146
rect -886 1103 -834 1112
rect -821 1103 -769 1112
rect -756 1103 -704 1112
rect -691 1146 -639 1155
rect -691 1112 -688 1146
rect -688 1112 -654 1146
rect -654 1112 -639 1146
rect -691 1103 -639 1112
rect -626 1146 -574 1155
rect -626 1112 -614 1146
rect -614 1112 -580 1146
rect -580 1112 -574 1146
rect -626 1103 -574 1112
rect -562 1146 -510 1155
rect -498 1146 -446 1155
rect -434 1146 -382 1155
rect -370 1146 -318 1155
rect -306 1146 -254 1155
rect -242 1146 -190 1155
rect -562 1112 -540 1146
rect -540 1112 -510 1146
rect -498 1112 -466 1146
rect -466 1112 -446 1146
rect -434 1112 -432 1146
rect -432 1112 -392 1146
rect -392 1112 -382 1146
rect -370 1112 -358 1146
rect -358 1112 -319 1146
rect -319 1112 -318 1146
rect -306 1112 -285 1146
rect -285 1112 -254 1146
rect -242 1112 -212 1146
rect -212 1112 -190 1146
rect -562 1103 -510 1112
rect -498 1103 -446 1112
rect -434 1103 -382 1112
rect -370 1103 -318 1112
rect -306 1103 -254 1112
rect -242 1103 -190 1112
rect -178 1146 -126 1155
rect -178 1112 -173 1146
rect -173 1112 -139 1146
rect -139 1112 -126 1146
rect -178 1103 -126 1112
rect -114 1146 -62 1155
rect -114 1112 -100 1146
rect -100 1112 -66 1146
rect -66 1112 -62 1146
rect -114 1103 -62 1112
rect -50 1146 2 1155
rect 14 1146 66 1155
rect 78 1146 130 1155
rect 142 1146 194 1155
rect 206 1146 258 1155
rect 270 1146 322 1155
rect -50 1112 -27 1146
rect -27 1112 2 1146
rect 14 1112 46 1146
rect 46 1112 66 1146
rect 78 1112 80 1146
rect 80 1112 119 1146
rect 119 1112 130 1146
rect 142 1112 153 1146
rect 153 1112 192 1146
rect 192 1112 194 1146
rect 206 1112 226 1146
rect 226 1112 258 1146
rect 270 1112 299 1146
rect 299 1112 322 1146
rect -50 1103 2 1112
rect 14 1103 66 1112
rect 78 1103 130 1112
rect 142 1103 194 1112
rect 206 1103 258 1112
rect 270 1103 322 1112
rect 334 1146 386 1155
rect 334 1112 338 1146
rect 338 1112 372 1146
rect 372 1112 386 1146
rect 334 1103 386 1112
rect 398 1146 450 1155
rect 398 1112 411 1146
rect 411 1112 445 1146
rect 445 1112 450 1146
rect 398 1103 450 1112
rect 462 1146 514 1155
rect 526 1146 578 1155
rect 590 1146 642 1155
rect 654 1146 706 1155
rect 462 1112 484 1146
rect 484 1112 514 1146
rect 526 1112 557 1146
rect 557 1112 578 1146
rect 590 1112 591 1146
rect 591 1112 630 1146
rect 630 1112 642 1146
rect 654 1112 664 1146
rect 664 1112 703 1146
rect 703 1112 706 1146
rect 462 1103 514 1112
rect 526 1103 578 1112
rect 590 1103 642 1112
rect 654 1103 706 1112
rect -886 1072 -834 1083
rect -821 1072 -769 1083
rect -756 1072 -704 1083
rect -886 1038 -876 1072
rect -876 1038 -836 1072
rect -836 1038 -834 1072
rect -821 1038 -802 1072
rect -802 1038 -769 1072
rect -756 1038 -728 1072
rect -728 1038 -704 1072
rect -886 1031 -834 1038
rect -821 1031 -769 1038
rect -756 1031 -704 1038
rect -691 1072 -639 1083
rect -691 1038 -688 1072
rect -688 1038 -654 1072
rect -654 1038 -639 1072
rect -691 1031 -639 1038
rect -626 1072 -574 1083
rect -626 1038 -614 1072
rect -614 1038 -580 1072
rect -580 1038 -574 1072
rect -626 1031 -574 1038
rect -562 1072 -510 1083
rect -498 1072 -446 1083
rect -434 1072 -382 1083
rect -370 1072 -318 1083
rect -306 1072 -254 1083
rect -242 1072 -190 1083
rect -562 1038 -540 1072
rect -540 1038 -510 1072
rect -498 1038 -466 1072
rect -466 1038 -446 1072
rect -434 1038 -432 1072
rect -432 1038 -392 1072
rect -392 1038 -382 1072
rect -370 1038 -358 1072
rect -358 1038 -319 1072
rect -319 1038 -318 1072
rect -306 1038 -285 1072
rect -285 1038 -254 1072
rect -242 1038 -212 1072
rect -212 1038 -190 1072
rect -562 1031 -510 1038
rect -498 1031 -446 1038
rect -434 1031 -382 1038
rect -370 1031 -318 1038
rect -306 1031 -254 1038
rect -242 1031 -190 1038
rect -178 1072 -126 1083
rect -178 1038 -173 1072
rect -173 1038 -139 1072
rect -139 1038 -126 1072
rect -178 1031 -126 1038
rect -114 1072 -62 1083
rect -114 1038 -100 1072
rect -100 1038 -66 1072
rect -66 1038 -62 1072
rect -114 1031 -62 1038
rect -50 1072 2 1083
rect 14 1072 66 1083
rect 78 1072 130 1083
rect 142 1072 194 1083
rect 206 1072 258 1083
rect 270 1072 322 1083
rect -50 1038 -27 1072
rect -27 1038 2 1072
rect 14 1038 46 1072
rect 46 1038 66 1072
rect 78 1038 80 1072
rect 80 1038 119 1072
rect 119 1038 130 1072
rect 142 1038 153 1072
rect 153 1038 192 1072
rect 192 1038 194 1072
rect 206 1038 226 1072
rect 226 1038 258 1072
rect 270 1038 299 1072
rect 299 1038 322 1072
rect -50 1031 2 1038
rect 14 1031 66 1038
rect 78 1031 130 1038
rect 142 1031 194 1038
rect 206 1031 258 1038
rect 270 1031 322 1038
rect 334 1072 386 1083
rect 334 1038 338 1072
rect 338 1038 372 1072
rect 372 1038 386 1072
rect 334 1031 386 1038
rect 398 1072 450 1083
rect 398 1038 411 1072
rect 411 1038 445 1072
rect 445 1038 450 1072
rect 398 1031 450 1038
rect 462 1072 514 1083
rect 526 1072 578 1083
rect 590 1072 642 1083
rect 654 1072 706 1083
rect 462 1038 484 1072
rect 484 1038 514 1072
rect 526 1038 557 1072
rect 557 1038 578 1072
rect 590 1038 591 1072
rect 591 1038 630 1072
rect 630 1038 642 1072
rect 654 1038 664 1072
rect 664 1038 703 1072
rect 703 1038 706 1072
rect 462 1031 514 1038
rect 526 1031 578 1038
rect 590 1031 642 1038
rect 654 1031 706 1038
rect -886 998 -834 1011
rect -821 998 -769 1011
rect -756 998 -704 1011
rect -886 964 -876 998
rect -876 964 -836 998
rect -836 964 -834 998
rect -821 964 -802 998
rect -802 964 -769 998
rect -756 964 -728 998
rect -728 964 -704 998
rect -886 959 -834 964
rect -821 959 -769 964
rect -756 959 -704 964
rect -691 998 -639 1011
rect -691 964 -688 998
rect -688 964 -654 998
rect -654 964 -639 998
rect -691 959 -639 964
rect -626 998 -574 1011
rect -626 964 -614 998
rect -614 964 -580 998
rect -580 964 -574 998
rect -626 959 -574 964
rect -562 998 -510 1011
rect -498 998 -446 1011
rect -434 998 -382 1011
rect -370 998 -318 1011
rect -306 998 -254 1011
rect -242 998 -190 1011
rect -562 964 -540 998
rect -540 964 -510 998
rect -498 964 -466 998
rect -466 964 -446 998
rect -434 964 -432 998
rect -432 964 -392 998
rect -392 964 -382 998
rect -370 964 -358 998
rect -358 964 -319 998
rect -319 964 -318 998
rect -306 964 -285 998
rect -285 964 -254 998
rect -242 964 -212 998
rect -212 964 -190 998
rect -562 959 -510 964
rect -498 959 -446 964
rect -434 959 -382 964
rect -370 959 -318 964
rect -306 959 -254 964
rect -242 959 -190 964
rect -178 998 -126 1011
rect -178 964 -173 998
rect -173 964 -139 998
rect -139 964 -126 998
rect -178 959 -126 964
rect -114 998 -62 1011
rect -114 964 -100 998
rect -100 964 -66 998
rect -66 964 -62 998
rect -114 959 -62 964
rect -50 998 2 1011
rect 14 998 66 1011
rect 78 998 130 1011
rect 142 998 194 1011
rect 206 998 258 1011
rect 270 998 322 1011
rect -50 964 -27 998
rect -27 964 2 998
rect 14 964 46 998
rect 46 964 66 998
rect 78 964 80 998
rect 80 964 119 998
rect 119 964 130 998
rect 142 964 153 998
rect 153 964 192 998
rect 192 964 194 998
rect 206 964 226 998
rect 226 964 258 998
rect 270 964 299 998
rect 299 964 322 998
rect -50 959 2 964
rect 14 959 66 964
rect 78 959 130 964
rect 142 959 194 964
rect 206 959 258 964
rect 270 959 322 964
rect 334 998 386 1011
rect 334 964 338 998
rect 338 964 372 998
rect 372 964 386 998
rect 334 959 386 964
rect 398 998 450 1011
rect 398 964 411 998
rect 411 964 445 998
rect 445 964 450 998
rect 398 959 450 964
rect 462 998 514 1011
rect 526 998 578 1011
rect 590 998 642 1011
rect 654 998 706 1011
rect 462 964 484 998
rect 484 964 514 998
rect 526 964 557 998
rect 557 964 578 998
rect 590 964 591 998
rect 591 964 630 998
rect 630 964 642 998
rect 654 964 664 998
rect 664 964 703 998
rect 703 964 706 998
rect 462 959 514 964
rect 526 959 578 964
rect 590 959 642 964
rect 654 959 706 964
rect 18784 946 18964 1126
rect 24755 1068 24807 1120
rect 24819 1068 24871 1120
rect 23954 989 24006 1041
rect 24019 989 24071 1041
rect -886 924 -834 939
rect -821 924 -769 939
rect -756 924 -704 939
rect -886 890 -876 924
rect -876 890 -836 924
rect -836 890 -834 924
rect -821 890 -802 924
rect -802 890 -769 924
rect -756 890 -728 924
rect -728 890 -704 924
rect -886 887 -834 890
rect -821 887 -769 890
rect -756 887 -704 890
rect -691 924 -639 939
rect -691 890 -688 924
rect -688 890 -654 924
rect -654 890 -639 924
rect -691 887 -639 890
rect -626 924 -574 939
rect -626 890 -614 924
rect -614 890 -580 924
rect -580 890 -574 924
rect -626 887 -574 890
rect -562 924 -510 939
rect -498 924 -446 939
rect -434 924 -382 939
rect -370 924 -318 939
rect -306 924 -254 939
rect -242 924 -190 939
rect -562 890 -540 924
rect -540 890 -510 924
rect -498 890 -466 924
rect -466 890 -446 924
rect -434 890 -432 924
rect -432 890 -392 924
rect -392 890 -382 924
rect -370 890 -358 924
rect -358 890 -319 924
rect -319 890 -318 924
rect -306 890 -285 924
rect -285 890 -254 924
rect -242 890 -212 924
rect -212 890 -190 924
rect -562 887 -510 890
rect -498 887 -446 890
rect -434 887 -382 890
rect -370 887 -318 890
rect -306 887 -254 890
rect -242 887 -190 890
rect -178 924 -126 939
rect -178 890 -173 924
rect -173 890 -139 924
rect -139 890 -126 924
rect -178 887 -126 890
rect -114 924 -62 939
rect -114 890 -100 924
rect -100 890 -66 924
rect -66 890 -62 924
rect -114 887 -62 890
rect -50 924 2 939
rect 14 924 66 939
rect 78 924 130 939
rect 142 924 194 939
rect 206 924 258 939
rect 270 924 322 939
rect -50 890 -27 924
rect -27 890 2 924
rect 14 890 46 924
rect 46 890 66 924
rect 78 890 80 924
rect 80 890 119 924
rect 119 890 130 924
rect 142 890 153 924
rect 153 890 192 924
rect 192 890 194 924
rect 206 890 226 924
rect 226 890 258 924
rect 270 890 299 924
rect 299 890 322 924
rect -50 887 2 890
rect 14 887 66 890
rect 78 887 130 890
rect 142 887 194 890
rect 206 887 258 890
rect 270 887 322 890
rect 334 924 386 939
rect 334 890 338 924
rect 338 890 372 924
rect 372 890 386 924
rect 334 887 386 890
rect 398 924 450 939
rect 398 890 411 924
rect 411 890 445 924
rect 445 890 450 924
rect 398 887 450 890
rect 462 924 514 939
rect 526 924 578 939
rect 590 924 642 939
rect 654 924 706 939
rect 462 890 484 924
rect 484 890 514 924
rect 526 890 557 924
rect 557 890 578 924
rect 590 890 591 924
rect 591 890 630 924
rect 630 890 642 924
rect 654 890 664 924
rect 664 890 703 924
rect 703 890 706 924
rect 462 887 514 890
rect 526 887 578 890
rect 590 887 642 890
rect 654 887 706 890
rect -886 850 -834 867
rect -821 850 -769 867
rect -756 850 -704 867
rect -886 816 -876 850
rect -876 816 -836 850
rect -836 816 -834 850
rect -821 816 -802 850
rect -802 816 -769 850
rect -756 816 -728 850
rect -728 816 -704 850
rect -886 815 -834 816
rect -821 815 -769 816
rect -756 815 -704 816
rect -691 850 -639 867
rect -691 816 -688 850
rect -688 816 -654 850
rect -654 816 -639 850
rect -691 815 -639 816
rect -626 850 -574 867
rect -626 816 -614 850
rect -614 816 -580 850
rect -580 816 -574 850
rect -626 815 -574 816
rect -562 850 -510 867
rect -498 850 -446 867
rect -434 850 -382 867
rect -370 850 -318 867
rect -306 850 -254 867
rect -242 850 -190 867
rect -562 816 -540 850
rect -540 816 -510 850
rect -498 816 -466 850
rect -466 816 -446 850
rect -434 816 -432 850
rect -432 816 -392 850
rect -392 816 -382 850
rect -370 816 -358 850
rect -358 816 -319 850
rect -319 816 -318 850
rect -306 816 -285 850
rect -285 816 -254 850
rect -242 816 -212 850
rect -212 816 -190 850
rect -562 815 -510 816
rect -498 815 -446 816
rect -434 815 -382 816
rect -370 815 -318 816
rect -306 815 -254 816
rect -242 815 -190 816
rect -178 850 -126 867
rect -178 816 -173 850
rect -173 816 -139 850
rect -139 816 -126 850
rect -178 815 -126 816
rect -114 850 -62 867
rect -114 816 -100 850
rect -100 816 -66 850
rect -66 816 -62 850
rect -114 815 -62 816
rect -50 850 2 867
rect 14 850 66 867
rect 78 850 130 867
rect 142 850 194 867
rect 206 850 258 867
rect 270 850 322 867
rect -50 816 -27 850
rect -27 816 2 850
rect 14 816 46 850
rect 46 816 66 850
rect 78 816 80 850
rect 80 816 119 850
rect 119 816 130 850
rect 142 816 153 850
rect 153 816 192 850
rect 192 816 194 850
rect 206 816 226 850
rect 226 816 258 850
rect 270 816 299 850
rect 299 816 322 850
rect -50 815 2 816
rect 14 815 66 816
rect 78 815 130 816
rect 142 815 194 816
rect 206 815 258 816
rect 270 815 322 816
rect 334 850 386 867
rect 334 816 338 850
rect 338 816 372 850
rect 372 816 386 850
rect 334 815 386 816
rect 398 850 450 867
rect 398 816 411 850
rect 411 816 445 850
rect 445 816 450 850
rect 398 815 450 816
rect 462 850 514 867
rect 526 850 578 867
rect 590 850 642 867
rect 654 850 706 867
rect 462 816 484 850
rect 484 816 514 850
rect 526 816 557 850
rect 557 816 578 850
rect 590 816 591 850
rect 591 816 630 850
rect 630 816 642 850
rect 654 816 664 850
rect 664 816 703 850
rect 703 816 706 850
rect 462 815 514 816
rect 526 815 578 816
rect 590 815 642 816
rect 654 815 706 816
rect 24057 934 24109 943
rect 24057 900 24090 934
rect 24090 900 24109 934
rect 24057 891 24109 900
rect 24121 934 24173 943
rect 24121 900 24128 934
rect 24128 900 24162 934
rect 24162 900 24173 934
rect 24121 891 24173 900
rect 24343 934 24395 943
rect 24343 900 24347 934
rect 24347 900 24381 934
rect 24381 900 24395 934
rect 24343 891 24395 900
rect 24407 934 24459 943
rect 24407 900 24419 934
rect 24419 900 24453 934
rect 24453 900 24459 934
rect 24407 891 24459 900
rect 24624 934 24676 943
rect 24624 900 24630 934
rect 24630 900 24664 934
rect 24664 900 24676 934
rect 24624 891 24676 900
rect 24688 934 24740 943
rect 24688 900 24702 934
rect 24702 900 24736 934
rect 24736 900 24740 934
rect 24688 891 24740 900
rect 24931 927 24983 961
rect 24931 909 24937 927
rect 24937 909 24971 927
rect 24971 909 24983 927
rect 24995 927 25047 961
rect 24995 909 25009 927
rect 25009 909 25043 927
rect 25043 909 25047 927
rect 25101 893 25153 899
rect 25101 859 25107 893
rect 25107 859 25141 893
rect 25141 859 25153 893
rect 25101 847 25153 859
rect 25165 893 25217 899
rect 25165 859 25179 893
rect 25179 859 25213 893
rect 25213 859 25217 893
rect 25165 847 25217 859
rect 25645 859 25697 911
rect 25645 795 25697 847
rect 24833 689 24885 741
rect 24897 689 24949 741
rect 24501 615 24507 649
rect 24507 615 24541 649
rect 24541 615 24553 649
rect 24501 597 24553 615
rect 23283 494 23335 546
rect 23347 494 23399 546
rect 24501 511 24553 563
rect -730 167 -678 219
rect -247 177 -195 229
rect -183 177 -131 229
rect -730 103 -678 155
rect 19413 129 19465 181
rect 19477 129 19529 181
rect 13237 -65 13289 -13
rect 13304 -65 13356 -13
rect 13371 -65 13423 -13
rect 13438 -65 13490 -13
rect 13505 -65 13557 -13
rect 13572 -65 13624 -13
rect 13639 -65 13691 -13
rect 13705 -65 13757 -13
rect 13771 -65 13823 -13
rect 13237 -169 13289 -117
rect 13304 -169 13356 -117
rect 13371 -169 13423 -117
rect 13438 -169 13490 -117
rect 13505 -169 13557 -117
rect 13572 -169 13624 -117
rect 13639 -169 13691 -117
rect 13705 -169 13757 -117
rect 13771 -169 13823 -117
rect 641 -4413 693 -4361
rect 707 -4413 759 -4361
<< metal2 >>
rect 1357 22407 2335 22413
rect 1409 22355 1513 22407
rect 1565 22355 2335 22407
rect 1357 22343 2335 22355
rect 1409 22291 1513 22343
rect 1565 22291 2335 22343
rect 1357 22285 2335 22291
tri 2120 22251 2154 22285 ne
rect 2154 22251 2335 22285
rect 1435 22245 1487 22251
tri 2154 22201 2204 22251 ne
rect 1435 22181 1487 22193
rect 1435 22117 1487 22129
tri 1404 22009 1435 22040 se
rect 1435 22009 1487 22065
rect 1176 21957 1487 22009
tri 1157 21251 1176 21270 se
rect 1176 21251 1228 21957
tri 1228 21926 1259 21957 nw
rect 1279 21907 2164 21913
rect 1331 21855 1591 21907
rect 1643 21855 2164 21907
rect 1279 21843 2164 21855
rect 1331 21791 1591 21843
rect 1643 21791 2164 21843
rect 1279 21779 2164 21791
rect 1331 21727 1591 21779
rect 1643 21727 2164 21779
rect 1279 21721 2164 21727
tri 2073 21682 2112 21721 ne
rect 1279 21583 2072 21589
rect 1331 21531 1591 21583
rect 1643 21531 2072 21583
rect 1279 21519 2072 21531
rect 1331 21467 1591 21519
rect 1643 21467 2072 21519
rect 1279 21455 2072 21467
rect 1331 21403 1591 21455
rect 1643 21403 2072 21455
rect 1279 21397 2072 21403
tri 1984 21361 2020 21397 ne
tri 1151 21245 1157 21251 se
rect 1157 21245 1228 21251
tri 1145 21239 1151 21245 se
rect 1151 21239 1228 21245
rect 449 21187 1228 21239
rect 1435 21245 1487 21251
rect 449 21181 527 21187
tri 527 21181 533 21187 nw
rect 1435 21181 1487 21193
rect 449 21172 518 21181
tri 518 21172 527 21181 nw
tri 422 15847 449 15874 se
rect 449 15847 501 21172
tri 501 21155 518 21172 nw
tri 1418 21155 1435 21172 se
tri 1405 21142 1418 21155 se
rect 1418 21142 1435 21155
rect 295 15832 501 15847
rect 295 15795 464 15832
tri 464 15795 501 15832 nw
rect 539 21129 1435 21142
rect 539 21117 1487 21129
rect 539 21090 1435 21117
rect 539 21065 598 21090
tri 598 21065 623 21090 nw
tri 1404 21065 1429 21090 ne
rect 1429 21065 1435 21090
rect 539 21059 592 21065
tri 592 21059 598 21065 nw
tri 1429 21059 1435 21065 ne
rect 1435 21059 1487 21065
rect 295 9466 347 15795
rect 539 15757 591 21059
tri 591 21058 592 21059 nw
rect 379 15705 591 15757
rect 379 10150 431 15705
rect 2020 14640 2072 21397
rect 2020 14565 2072 14588
rect 2020 14507 2072 14513
rect 2112 14640 2164 21721
rect 2204 14916 2335 22251
rect 2112 14565 2164 14588
rect 2112 14507 2164 14513
rect 1341 14302 1393 14308
rect 1341 14227 1393 14250
rect 1341 10756 1393 14175
rect 1341 10689 1393 10704
rect 379 10098 1215 10150
rect 1163 10074 1215 10098
rect 1163 10010 1215 10022
rect 1163 9952 1215 9958
rect 295 9460 1215 9466
rect 295 9414 1163 9460
rect 1163 9396 1215 9408
rect 1163 9338 1215 9344
rect 1341 9287 1393 10637
rect 1433 14300 1485 14306
rect 1433 14225 1485 14248
rect 1433 9697 1485 14173
rect 2159 12060 2211 12224
rect 2374 12087 2471 12139
tri 2392 12071 2408 12087 ne
rect 2408 12071 2471 12087
tri 2211 12060 2222 12071 sw
tri 2408 12060 2419 12071 ne
rect 2159 12059 2222 12060
tri 2222 12059 2223 12060 sw
rect 2159 12039 2223 12059
tri 2159 12027 2171 12039 ne
rect 1678 10756 1730 10762
rect 1678 10689 1730 10704
rect 1678 10505 1730 10637
rect 1678 10435 1730 10453
rect 1678 10364 1730 10383
rect 1678 10306 1730 10312
rect 1433 9627 1485 9645
rect 1433 9556 1485 9575
rect 1433 9298 1485 9504
rect 2171 10074 2223 12039
rect 2171 10010 2223 10022
tri 1433 9288 1443 9298 ne
rect 1443 9288 1485 9298
tri 1393 9287 1394 9288 sw
tri 1443 9287 1444 9288 ne
rect 1444 9287 1485 9288
rect 1341 9274 1394 9287
tri 1341 9237 1378 9274 ne
rect 1378 9249 1394 9274
tri 1394 9249 1432 9287 sw
tri 1444 9249 1482 9287 ne
rect 1482 9249 1485 9287
tri 1485 9249 1547 9311 sw
rect 1378 9246 1432 9249
tri 1432 9246 1435 9249 sw
tri 1482 9246 1485 9249 ne
rect 1485 9246 1547 9249
rect 1378 9237 1435 9246
tri 1435 9237 1444 9246 sw
tri 1485 9237 1494 9246 ne
rect 1494 9237 1547 9246
tri 1378 9222 1393 9237 ne
rect 1393 9222 1444 9237
tri 1393 9171 1444 9222 ne
tri 1444 9221 1460 9237 sw
tri 1494 9221 1510 9237 ne
rect 1510 9221 1547 9237
rect 1444 9184 1460 9221
tri 1460 9184 1497 9221 sw
tri 1510 9184 1547 9221 ne
tri 1547 9184 1612 9249 sw
rect 2171 9184 2223 9958
rect 2337 9514 2389 11575
rect 2419 10541 2471 12071
rect 2419 10477 2471 10489
rect 2419 9870 2471 10425
rect 2419 9806 2471 9818
rect 2419 9663 2471 9754
rect 2337 9450 2389 9462
tri 2223 9184 2231 9192 sw
rect 1444 9171 1497 9184
tri 1497 9171 1510 9184 sw
tri 1547 9171 1560 9184 ne
rect 1560 9171 1612 9184
tri 1444 9105 1510 9171 ne
tri 1510 9155 1526 9171 sw
tri 1560 9155 1576 9171 ne
rect 1576 9155 1612 9171
rect 1510 9119 1526 9155
tri 1526 9119 1562 9155 sw
tri 1576 9119 1612 9155 ne
tri 1612 9119 1677 9184 sw
rect 2171 9178 2231 9184
tri 2171 9174 2175 9178 ne
rect 2175 9174 2231 9178
tri 2231 9174 2241 9184 sw
tri 2175 9126 2223 9174 ne
rect 2223 9126 2241 9174
tri 2223 9119 2230 9126 ne
rect 2230 9119 2241 9126
tri 2241 9119 2296 9174 sw
rect 1510 9105 1562 9119
tri 1562 9105 1576 9119 sw
tri 1612 9105 1626 9119 ne
rect 1626 9105 2166 9119
tri 1510 9039 1576 9105 ne
tri 1576 9089 1592 9105 sw
tri 1626 9089 1642 9105 ne
rect 1642 9089 2166 9105
rect 1576 9069 1592 9089
tri 1592 9069 1612 9089 sw
tri 1642 9069 1662 9089 ne
rect 1662 9069 2166 9089
rect 1576 9063 1612 9069
tri 1612 9063 1618 9069 sw
tri 2136 9063 2142 9069 ne
rect 2142 9063 2166 9069
tri 2166 9063 2222 9119 sw
tri 2230 9108 2241 9119 ne
rect 2241 9108 2296 9119
tri 2296 9108 2307 9119 sw
tri 2241 9094 2255 9108 ne
rect 1576 9039 1618 9063
tri 1618 9039 1642 9063 sw
tri 2142 9039 2166 9063 ne
rect 2166 9039 2222 9063
tri 1576 9008 1607 9039 ne
rect 1607 9035 2099 9039
tri 2099 9035 2103 9039 sw
tri 2166 9035 2170 9039 ne
rect 1607 9008 2103 9035
tri 2103 9008 2130 9035 sw
tri 1607 8997 1618 9008 ne
rect 1618 8997 2130 9008
tri 2044 8963 2078 8997 ne
tri 2009 6388 2078 6457 se
rect 2078 6439 2130 8997
rect 2078 6388 2079 6439
tri 2079 6388 2130 6439 nw
tri 2008 6387 2009 6388 se
rect 2009 6387 2078 6388
tri 2078 6387 2079 6388 nw
tri 2002 6381 2008 6387 se
rect 2008 6381 2072 6387
tri 2072 6381 2078 6387 nw
tri 1983 6281 2002 6300 se
rect 2002 6281 2054 6381
tri 2054 6363 2072 6381 nw
tri 2159 6363 2170 6374 se
rect 2170 6363 2222 9039
tri 2132 6336 2159 6363 se
rect 2159 6336 2222 6363
tri 2129 6333 2132 6336 se
rect 2132 6333 2222 6336
rect 2094 6281 2100 6333
rect 2152 6281 2164 6333
rect 2216 6281 2222 6333
tri 1961 6259 1983 6281 se
rect 1983 6259 2054 6281
rect 1926 6207 1932 6259
rect 1984 6207 1996 6259
rect 2048 6207 2054 6259
rect 2255 5988 2307 9108
rect 2255 5924 2307 5936
rect 2255 5866 2307 5872
rect 2337 5918 2389 9398
rect 15679 8055 15984 8064
rect 8094 7899 8103 7955
rect 8159 7899 8193 7955
rect 8249 7899 8283 7955
rect 8339 7899 8372 7955
rect 8428 7899 8461 7955
rect 8517 7899 8526 7955
rect 8094 7875 8526 7899
rect 8094 7819 8103 7875
rect 8159 7819 8193 7875
rect 8249 7819 8283 7875
rect 8339 7819 8372 7875
rect 8428 7819 8461 7875
rect 8517 7819 8526 7875
tri 7144 7778 7185 7819 se
rect 7185 7778 7392 7819
rect 6575 7769 7392 7778
rect 6711 7666 7392 7769
rect 8094 7795 8526 7819
rect 8094 7739 8103 7795
rect 8159 7739 8193 7795
rect 8249 7739 8283 7795
rect 8339 7739 8372 7795
rect 8428 7739 8461 7795
rect 8517 7739 8526 7795
rect 12741 7899 12750 7955
rect 12806 7899 12840 7955
rect 12896 7899 12930 7955
rect 12986 7899 13019 7955
rect 13075 7899 13108 7955
rect 13164 7899 13378 7955
rect 12741 7875 13378 7899
rect 12741 7819 12750 7875
rect 12806 7819 12840 7875
rect 12896 7819 12930 7875
rect 12986 7819 13019 7875
rect 13075 7819 13108 7875
rect 13164 7819 13378 7875
rect 12741 7795 13378 7819
rect 12741 7739 12750 7795
rect 12806 7739 12840 7795
rect 12896 7739 12930 7795
rect 12986 7739 13019 7795
rect 13075 7739 13108 7795
rect 13164 7739 13378 7795
rect 14270 7899 14279 7955
rect 14335 7899 14367 7955
rect 14423 7899 14455 7955
rect 14511 7899 14543 7955
rect 14599 7899 14630 7955
rect 14686 7899 14695 7955
rect 14270 7875 14695 7899
rect 14270 7819 14279 7875
rect 14335 7819 14367 7875
rect 14423 7819 14455 7875
rect 14511 7819 14543 7875
rect 14599 7819 14630 7875
rect 14686 7819 14695 7875
rect 14270 7795 14695 7819
rect 14270 7739 14279 7795
rect 14335 7739 14367 7795
rect 14423 7739 14455 7795
rect 14511 7739 14543 7795
rect 14599 7739 14630 7795
rect 14686 7739 14695 7795
rect 15679 7839 15846 8055
rect 15982 7839 15984 8055
rect 15679 7830 15984 7839
rect 15679 7739 15757 7830
tri 15757 7739 15848 7830 nw
tri 9144 7682 9171 7709 se
rect 9171 7682 9301 7685
rect 6711 7663 7389 7666
tri 7389 7663 7392 7666 nw
tri 8715 7663 8734 7682 se
rect 8734 7663 9301 7682
rect 12741 7663 13378 7739
rect 15679 7663 15681 7739
tri 15681 7663 15757 7739 nw
rect 6711 7659 7385 7663
tri 7385 7659 7389 7663 nw
tri 8711 7659 8715 7663 se
rect 8715 7659 9301 7663
tri 15679 7661 15681 7663 nw
rect 6711 7553 7270 7659
rect 6575 7544 7270 7553
tri 7270 7544 7385 7659 nw
tri 8698 7646 8711 7659 se
rect 8711 7657 9301 7659
rect 8711 7646 9290 7657
tri 9290 7646 9301 7657 nw
rect 8698 7616 9260 7646
tri 9260 7616 9290 7646 nw
rect 8698 6030 8748 7616
tri 8748 7587 8777 7616 nw
tri 13536 7547 13563 7574 se
rect 13563 7547 13693 7659
tri 13111 7523 13135 7547 se
rect 13135 7539 13693 7547
rect 13135 7523 13677 7539
tri 13677 7523 13693 7539 nw
rect 13111 7481 13635 7523
tri 13635 7481 13677 7523 nw
tri 8748 6030 8752 6034 sw
tri 8661 5993 8698 6030 se
rect 8698 5993 8752 6030
tri 8752 5993 8789 6030 sw
rect 8661 5941 8667 5993
rect 8719 5941 8731 5993
rect 8783 5941 8789 5993
tri 13108 5941 13111 5944 se
rect 13111 5941 13161 7481
tri 13161 7464 13178 7481 nw
tri 25223 6342 25269 6388 se
rect 25269 6342 25526 6388
rect 25223 6336 25526 6342
rect 25578 6336 25590 6388
rect 25642 6336 25648 6388
rect 25223 6311 25325 6336
tri 25325 6311 25350 6336 nw
rect 25063 6241 25069 6293
rect 25121 6241 25133 6293
rect 25185 6241 25191 6293
tri 25063 6209 25095 6241 ne
tri 13085 5918 13108 5941 se
rect 13108 5918 13161 5941
tri 13161 5918 13185 5942 sw
rect 2337 5866 2359 5918
rect 2411 5866 2423 5918
rect 2475 5866 2481 5918
rect 13058 5866 13064 5918
rect 13116 5866 13128 5918
rect 13180 5866 13186 5918
rect -901 5778 8102 5834
rect 8158 5778 8192 5834
rect 8248 5778 8282 5834
rect 8338 5778 8371 5834
rect 8427 5778 8460 5834
rect 8516 5778 14275 5834
rect 14331 5778 14365 5834
rect 14421 5778 14455 5834
rect 14511 5778 14544 5834
rect 14600 5778 14633 5834
rect 14689 5778 14698 5834
rect -901 5754 14698 5778
rect -901 5698 8102 5754
rect 8158 5698 8192 5754
rect 8248 5698 8282 5754
rect 8338 5698 8371 5754
rect 8427 5698 8460 5754
rect 8516 5698 14275 5754
rect 14331 5698 14365 5754
rect 14421 5698 14455 5754
rect 14511 5698 14544 5754
rect 14600 5698 14633 5754
rect 14689 5698 14698 5754
rect 15841 5728 17068 5737
rect -901 4951 -781 5698
tri -781 5663 -746 5698 nw
rect 15897 5672 15931 5728
rect 15987 5681 17068 5728
rect 17124 5681 17151 5737
rect 17207 5681 17234 5737
rect 17290 5681 17299 5737
rect 15987 5672 17299 5681
tri -917 3145 -900 3162 se
rect -900 3145 -781 4951
tri -948 3114 -917 3145 se
rect -917 3114 -781 3145
tri -949 3113 -948 3114 se
rect -948 3113 -781 3114
tri -968 3094 -949 3113 se
rect -949 3094 -781 3113
rect -968 3092 -781 3094
rect -968 3040 -962 3092
rect -910 3040 -877 3092
rect -825 3040 -781 3092
rect -968 3012 -781 3040
rect -968 2960 -962 3012
rect -910 2960 -877 3012
rect -825 2960 -781 3012
rect -738 5662 13170 5663
rect -738 5631 13173 5662
rect -738 5575 12750 5631
rect 12806 5575 12840 5631
rect 12896 5575 12930 5631
rect 12986 5575 13019 5631
rect 13075 5575 13108 5631
rect 13164 5575 13173 5631
rect -738 5544 13173 5575
rect 15841 5603 17299 5672
rect 15897 5547 15931 5603
rect 15987 5595 17299 5603
rect 15987 5547 17068 5595
rect -738 5538 -571 5544
tri -571 5538 -565 5544 nw
rect 15841 5539 17068 5547
rect 17124 5539 17151 5595
rect 17207 5539 17234 5595
rect 17290 5539 17299 5595
rect 15841 5538 17299 5539
rect -738 5507 -602 5538
tri -602 5507 -571 5538 nw
rect -738 3166 -617 5507
tri -617 5492 -602 5507 nw
rect 11081 5476 11407 5507
rect 11081 5420 11090 5476
rect 11146 5420 11174 5476
rect 11230 5420 11258 5476
rect 11314 5420 11342 5476
rect 11398 5420 11407 5476
rect 11081 5389 11407 5420
rect 13752 5476 14078 5507
rect 13752 5420 13761 5476
rect 13817 5420 13845 5476
rect 13901 5420 13929 5476
rect 13985 5420 14013 5476
rect 14069 5420 14078 5476
rect 13752 5389 14078 5420
rect -220 3310 -101 5235
rect 7342 5149 7348 5201
rect 7400 5149 7412 5201
rect 7464 5149 7888 5201
rect 7940 5149 7952 5201
rect 8004 5149 8010 5201
rect -52 3510 69 4929
rect 3757 4287 4086 5051
tri 17213 4601 17285 4673 nw
tri 17870 4601 17942 4673 ne
rect 21074 4287 21403 5051
tri 22346 4635 22380 4669 ne
rect 22380 4421 22412 4669
tri 22412 4635 22446 4669 nw
tri 22380 4411 22390 4421 ne
rect 22390 4411 22412 4421
tri 22412 4411 22436 4435 sw
tri 22390 4405 22396 4411 ne
rect 22396 4405 23456 4411
tri 23456 4405 23462 4411 sw
tri 22396 4389 22412 4405 ne
rect 22412 4389 23462 4405
tri 22412 4379 22422 4389 ne
rect 22422 4379 23462 4389
tri 23442 4359 23462 4379 ne
tri 23462 4359 23508 4405 sw
tri 23462 4313 23508 4359 ne
tri 23508 4313 23554 4359 sw
tri 23508 4287 23534 4313 ne
rect 23534 4287 23554 4313
tri 23554 4287 23580 4313 sw
tri 23534 4267 23554 4287 ne
rect 23554 4267 23580 4287
tri 23580 4267 23600 4287 sw
tri 23554 4261 23560 4267 ne
rect 23560 4261 24197 4267
tri 24197 4261 24203 4267 sw
tri 23560 4235 23586 4261 ne
rect 23586 4235 24203 4261
tri 24183 4215 24203 4235 ne
tri 24203 4215 24249 4261 sw
tri 24203 4207 24211 4215 ne
rect 24211 4207 24249 4215
tri 24249 4207 24257 4215 sw
rect 23422 4183 24099 4207
tri 24099 4183 24123 4207 sw
tri 24211 4183 24235 4207 ne
rect 24235 4183 24257 4207
tri 24257 4183 24281 4207 sw
rect 23422 4179 24123 4183
tri 24077 4138 24118 4179 ne
rect 24118 4138 24123 4179
rect 12187 4053 12233 4105
tri 12902 4079 12923 4100 se
rect 12930 4086 12968 4138
tri 24118 4133 24123 4138 ne
tri 24123 4133 24173 4183 sw
tri 24235 4169 24249 4183 ne
rect 24249 4169 24281 4183
tri 24281 4169 24295 4183 sw
tri 24249 4155 24263 4169 ne
tri 24123 4111 24145 4133 ne
rect 12902 4070 12975 4079
rect 12902 4014 12908 4070
rect 12964 4014 12975 4070
rect 12902 3986 12975 4014
rect 5392 3901 5401 3957
rect 5457 3901 5481 3957
rect 5537 3901 5546 3957
rect 12902 3930 12908 3986
rect 12964 3930 12975 3986
rect 12902 3917 12975 3930
rect 1094 3777 1146 3865
tri 1146 3777 1149 3780 sw
rect 1094 3747 1149 3777
tri 1149 3747 1179 3777 sw
tri 24004 3767 24014 3777 se
rect 24014 3767 24066 3865
tri 16855 3747 16867 3759 se
rect 16867 3747 16877 3759
rect 1094 3711 16877 3747
tri 16855 3703 16863 3711 ne
rect 16863 3703 16877 3711
rect 16933 3703 16957 3759
rect 17013 3703 17022 3759
rect 17442 3711 17451 3767
rect 17507 3711 17531 3767
rect 17587 3747 17596 3767
tri 17596 3747 17616 3767 sw
tri 23984 3747 24004 3767 se
rect 24004 3747 24066 3767
rect 17587 3711 24066 3747
tri 69 3510 78 3519 sw
rect 23224 3510 23230 3562
rect 23282 3510 23294 3562
rect 23346 3510 23352 3562
rect -52 3476 78 3510
tri 78 3476 112 3510 sw
rect -52 3431 112 3476
tri 112 3431 157 3476 sw
rect -52 3424 585 3431
tri 585 3424 592 3431 sw
rect 22871 3424 22877 3476
rect 22929 3424 22941 3476
rect 22993 3424 22999 3476
rect -52 3374 592 3424
tri 592 3374 642 3424 sw
rect -52 3343 642 3374
tri -52 3323 -32 3343 ne
rect -32 3323 642 3343
tri -101 3310 -88 3323 sw
tri -32 3310 -19 3323 ne
rect -19 3310 642 3323
rect -220 3286 -88 3310
tri -88 3286 -64 3310 sw
tri 222 3286 246 3310 ne
rect 246 3286 642 3310
rect -220 3257 -64 3286
tri -64 3257 -35 3286 sw
tri 246 3257 275 3286 ne
rect 275 3257 642 3286
rect -220 3205 -35 3257
tri -35 3205 17 3257 sw
tri 275 3205 327 3257 ne
rect 327 3205 642 3257
rect -220 3197 17 3205
tri 17 3197 25 3205 sw
tri 327 3197 335 3205 ne
rect 335 3197 642 3205
rect 12084 3267 12964 3276
rect 12140 3211 12908 3267
rect 12084 3204 12964 3211
rect -220 3181 25 3197
tri 25 3181 41 3197 sw
tri 335 3181 351 3197 ne
rect -220 3171 41 3181
tri 41 3171 51 3181 sw
tri -617 3166 -612 3171 sw
rect -220 3166 51 3171
tri 51 3166 56 3171 sw
rect -738 3145 -612 3166
tri -612 3145 -591 3166 sw
rect -220 3145 56 3166
tri 56 3145 77 3166 sw
rect -738 3114 -591 3145
tri -591 3114 -560 3145 sw
rect -220 3133 77 3145
tri -220 3114 -201 3133 ne
rect -201 3114 77 3133
tri 77 3114 108 3145 sw
rect -738 3113 -560 3114
tri -560 3113 -559 3114 sw
tri -201 3113 -200 3114 ne
rect -200 3113 108 3114
tri 108 3113 109 3114 sw
rect -738 3083 -559 3113
tri -559 3083 -529 3113 sw
tri -200 3083 -170 3113 ne
rect -170 3083 109 3113
tri 109 3083 139 3113 sw
rect -738 3056 -231 3083
tri -170 3076 -163 3083 ne
rect -163 3076 139 3083
tri 139 3076 146 3083 sw
tri -163 3062 -149 3076 ne
rect -149 3062 146 3076
tri -149 3061 -148 3062 ne
rect -148 3061 146 3062
tri -148 3060 -147 3061 ne
rect -738 3019 -617 3056
tri -738 3004 -723 3019 ne
rect -723 3004 -617 3019
rect -565 3004 -535 3056
rect -483 3004 -453 3056
rect -401 3004 -371 3056
rect -319 3004 -289 3056
rect -237 3004 -231 3056
tri -723 2986 -705 3004 ne
rect -705 2986 -231 3004
rect -147 3037 146 3061
rect -968 2932 -781 2960
rect -147 2985 -141 3037
rect -89 2985 -65 3037
rect -13 2985 11 3037
rect 63 2985 86 3037
rect 138 2985 146 3037
rect -147 2954 146 2985
rect 351 3037 642 3197
rect 10276 3142 10285 3198
rect 10341 3197 10367 3198
rect 10423 3197 10449 3198
rect 10505 3197 10530 3198
rect 10586 3197 10611 3198
rect 10667 3197 10692 3198
rect 10341 3145 10355 3197
rect 10679 3145 10692 3197
rect 10341 3142 10367 3145
rect 10423 3142 10449 3145
rect 10505 3142 10530 3145
rect 10586 3142 10611 3145
rect 10667 3142 10692 3145
rect 10748 3142 10757 3198
rect 10276 3113 10757 3142
rect 12084 3187 12141 3204
rect 12140 3166 12141 3187
tri 12141 3166 12179 3204 nw
tri 12869 3166 12907 3204 ne
rect 12907 3187 12964 3204
rect 12907 3166 12908 3187
tri 12140 3165 12141 3166 nw
tri 12907 3165 12908 3166 ne
rect 12084 3122 12140 3131
rect 12908 3122 12964 3131
rect 24145 3116 24173 4133
rect 24263 3211 24295 4169
tri 25066 3257 25095 3286 se
rect 25095 3259 25153 6241
tri 25153 6209 25185 6241 nw
rect 25095 3257 25151 3259
tri 25151 3257 25153 3259 nw
tri 24263 3205 24269 3211 ne
rect 24269 3205 24295 3211
tri 24295 3205 24315 3225 sw
rect 24513 3205 24519 3257
rect 24571 3205 24583 3257
rect 24635 3205 25099 3257
tri 25099 3205 25151 3257 nw
rect 25223 3223 25281 6311
tri 25281 6267 25325 6311 nw
rect 25416 5236 25468 5242
tri 25204 3205 25222 3223 se
rect 25222 3205 25281 3223
tri 24269 3182 24292 3205 ne
rect 24292 3182 24315 3205
tri 24315 3182 24338 3205 sw
tri 25181 3182 25204 3205 se
rect 25204 3182 25281 3205
tri 24292 3179 24295 3182 ne
rect 24295 3179 24338 3182
tri 24295 3166 24308 3179 ne
rect 24308 3166 24338 3179
tri 24338 3166 24354 3182 sw
tri 25165 3166 25181 3182 se
rect 25181 3166 25281 3182
tri 24308 3136 24338 3166 ne
rect 24338 3136 24354 3166
tri 24354 3136 24384 3166 sw
tri 24338 3132 24342 3136 ne
rect 24342 3132 24384 3136
tri 24384 3132 24388 3136 sw
tri 24145 3114 24147 3116 ne
rect 24147 3114 24173 3116
tri 24173 3114 24191 3132 sw
tri 24342 3114 24360 3132 ne
rect 24360 3114 24388 3132
tri 24388 3114 24406 3132 sw
rect 24520 3114 24526 3166
rect 24578 3114 24590 3166
rect 24642 3147 25281 3166
rect 24642 3114 25248 3147
tri 25248 3114 25281 3147 nw
rect 25325 5176 25377 5182
rect 25325 5096 25377 5124
rect 10276 3096 10286 3113
rect 10338 3096 10355 3113
rect 10407 3096 10423 3113
rect 10475 3096 10491 3113
rect 10543 3096 10559 3113
rect 10611 3096 10627 3113
rect 10679 3096 10695 3113
rect 10747 3096 10757 3113
tri 24147 3098 24163 3114 ne
rect 24163 3098 24191 3114
tri 24191 3098 24207 3114 sw
tri 24360 3098 24376 3114 ne
rect 24376 3098 24406 3114
tri 24406 3098 24422 3114 sw
rect 10276 3040 10285 3096
rect 10341 3061 10355 3096
rect 10679 3061 10692 3096
rect 10341 3040 10367 3061
rect 10423 3040 10449 3061
rect 10505 3040 10530 3061
rect 10586 3040 10611 3061
rect 10667 3040 10692 3061
rect 10748 3040 10757 3096
tri 24163 3088 24173 3098 ne
rect 24173 3088 24207 3098
tri 24173 3054 24207 3088 ne
tri 24207 3054 24251 3098 sw
tri 24376 3090 24384 3098 ne
rect 24384 3090 24422 3098
tri 24422 3090 24430 3098 sw
tri 24384 3054 24420 3090 ne
rect 24420 3054 24430 3090
tri 24430 3054 24466 3090 sw
tri 24207 3040 24221 3054 ne
rect 24221 3040 24251 3054
rect 351 2985 357 3037
rect 409 2985 433 3037
rect 485 2985 509 3037
rect 561 2985 584 3037
rect 636 2985 642 3037
tri 24221 3010 24251 3040 ne
tri 24251 3010 24295 3054 sw
tri 24420 3044 24430 3054 ne
rect 24430 3044 24466 3054
tri 24466 3044 24476 3054 sw
tri 24430 3010 24464 3044 ne
rect 24464 3010 24476 3044
tri 24476 3010 24510 3044 sw
tri 24251 3002 24259 3010 ne
rect 24259 3002 24369 3010
tri 24369 3002 24377 3010 sw
tri 24464 3002 24472 3010 ne
rect 24472 3002 24510 3010
tri 24510 3002 24518 3010 sw
rect 351 2956 642 2985
tri 24259 2982 24279 3002 ne
rect 24279 2982 24377 3002
tri 24349 2956 24375 2982 ne
rect 24375 2956 24377 2982
tri 24377 2956 24423 3002 sw
tri 24472 2998 24476 3002 ne
rect 24476 2998 24518 3002
tri 24518 2998 24522 3002 sw
tri 24476 2984 24490 2998 ne
tri 24375 2954 24377 2956 ne
rect 24377 2954 24423 2956
tri 24423 2954 24425 2956 sw
tri 24377 2934 24397 2954 ne
rect -968 2880 -962 2932
rect -910 2880 -877 2932
rect -825 2913 -781 2932
rect -825 2880 -819 2913
rect -968 2852 -819 2880
tri -819 2875 -781 2913 nw
rect -968 2800 -962 2852
rect -910 2800 -877 2852
rect -825 2800 -819 2852
rect 17360 2747 17806 2756
rect 17360 2745 17745 2747
rect 17360 2689 17365 2745
rect 17421 2691 17745 2745
rect 17801 2691 17806 2747
rect 17421 2689 17806 2691
rect 17360 2667 17806 2689
rect 17360 2665 17745 2667
rect 17360 2609 17365 2665
rect 17421 2611 17745 2665
rect 17801 2611 17806 2667
rect 17421 2609 17806 2611
rect 17360 2602 17806 2609
rect 17365 2600 17421 2602
rect 20734 2405 20743 2417
rect 20799 2405 20825 2417
rect 20881 2405 20907 2417
rect 20963 2405 20989 2417
rect 21045 2405 21071 2417
rect 21127 2405 21136 2417
rect 18842 2389 19116 2395
rect 18894 2337 18916 2389
rect 18968 2337 18990 2389
rect 19042 2337 19064 2389
rect 18842 2322 19116 2337
rect 18894 2319 18916 2322
rect 18968 2319 18990 2322
rect 19042 2319 19064 2322
rect 20734 2353 20742 2405
rect 20799 2361 20809 2405
rect 21062 2361 21071 2405
rect 20794 2353 20809 2361
rect 20861 2353 20876 2361
rect 20928 2353 20943 2361
rect 20995 2353 21010 2361
rect 21062 2353 21076 2361
rect 21128 2353 21136 2405
rect 20734 2337 21136 2353
rect 20734 2331 20743 2337
rect 20799 2331 20825 2337
rect 20881 2331 20907 2337
rect 20963 2331 20989 2337
rect 21045 2331 21071 2337
rect 21127 2331 21136 2337
rect 18839 2270 18842 2319
rect 18904 2270 18916 2319
rect 18839 2263 18848 2270
rect 18904 2263 18936 2270
rect 18992 2263 19024 2270
rect 19080 2263 19112 2270
rect 19168 2263 19177 2319
rect 18839 2255 19177 2263
rect 18839 2203 18842 2255
rect 18894 2203 18916 2255
rect 18968 2203 18990 2255
rect 19042 2203 19064 2255
rect 19116 2203 19177 2255
rect 18839 2193 19177 2203
rect 18839 2187 18848 2193
rect 18904 2187 18936 2193
rect 18992 2187 19024 2193
rect 19080 2187 19112 2193
rect 18839 2137 18842 2187
rect 18904 2137 18916 2187
rect 19168 2137 19177 2193
rect 20734 2279 20742 2331
rect 20799 2281 20809 2331
rect 21062 2281 21071 2331
rect 20794 2279 20809 2281
rect 20861 2279 20876 2281
rect 20928 2279 20943 2281
rect 20995 2279 21010 2281
rect 21062 2279 21076 2281
rect 21128 2279 21136 2331
rect 20734 2257 21136 2279
rect 20734 2205 20742 2257
rect 20799 2205 20809 2257
rect 21062 2205 21071 2257
rect 21128 2205 21136 2257
rect 20734 2201 20743 2205
rect 20799 2201 20825 2205
rect 20881 2201 20907 2205
rect 20963 2201 20989 2205
rect 21045 2201 21071 2205
rect 21127 2201 21136 2205
rect 20734 2183 21136 2201
rect 18894 2135 18916 2137
rect 18968 2135 18990 2137
rect 19042 2135 19064 2137
rect 18842 2119 19116 2135
rect 18894 2067 18916 2119
rect 18968 2067 18990 2119
rect 19042 2067 19064 2119
rect 18842 2061 19116 2067
rect 20734 2131 20742 2183
rect 20794 2177 20809 2183
rect 20861 2177 20876 2183
rect 20928 2177 20943 2183
rect 20995 2177 21010 2183
rect 21062 2177 21076 2183
rect 20799 2131 20809 2177
rect 21062 2131 21071 2177
rect 21128 2131 21136 2183
rect 20734 2121 20743 2131
rect 20799 2121 20825 2131
rect 20881 2121 20907 2131
rect 20963 2121 20989 2131
rect 21045 2121 21071 2131
rect 21127 2121 21136 2131
rect 20734 2109 21136 2121
rect 20734 2057 20742 2109
rect 20794 2097 20809 2109
rect 20861 2097 20876 2109
rect 20928 2097 20943 2109
rect 20995 2097 21010 2109
rect 21062 2097 21076 2109
rect 20799 2057 20809 2097
rect 21062 2057 21071 2097
rect 21128 2057 21136 2109
rect 20734 2041 20743 2057
rect 20799 2041 20825 2057
rect 20881 2041 20907 2057
rect 20963 2041 20989 2057
rect 21045 2041 21071 2057
rect 21127 2041 21136 2057
rect 1307 1872 1347 1924
rect 10348 1613 10354 1665
rect 10413 1613 10421 1665
rect 10473 1613 10480 1665
rect 10539 1613 10545 1665
rect 10348 1609 10357 1613
rect 10413 1609 10480 1613
rect 10536 1609 10545 1613
rect 10348 1573 10545 1609
rect 10348 1521 10354 1573
rect 10406 1563 10421 1573
rect 10413 1521 10421 1563
rect 10473 1563 10487 1573
rect 10473 1521 10480 1563
rect 10539 1521 10545 1573
rect 10348 1507 10357 1521
rect 10413 1507 10480 1521
rect 10536 1507 10545 1521
rect 24397 1576 24425 2954
tri 24425 1576 24449 1600 sw
rect 24397 1570 24449 1576
rect 24397 1505 24449 1518
rect 12084 1460 12140 1469
rect 24397 1447 24449 1453
rect 24397 1445 24447 1447
tri 24447 1445 24449 1447 nw
rect 12084 1380 12140 1404
tri 24376 1402 24397 1423 se
rect 24397 1402 24425 1445
tri 24425 1423 24447 1445 nw
rect 21019 1383 21042 1402
tri 24357 1383 24376 1402 se
rect 24376 1401 24425 1402
rect 24376 1383 24397 1401
tri 24347 1373 24357 1383 se
rect 24357 1373 24397 1383
tri 24397 1373 24425 1401 nw
tri 24341 1367 24347 1373 se
rect 24347 1367 24391 1373
tri 24391 1367 24397 1373 nw
tri 24335 1361 24341 1367 se
rect 24341 1361 24385 1367
tri 24385 1361 24391 1367 nw
tri 24299 1325 24335 1361 se
rect 24335 1325 24347 1361
rect 12084 1315 12140 1324
rect -892 1299 712 1301
rect -892 1247 -886 1299
rect -834 1247 -821 1299
rect -769 1247 -756 1299
rect -704 1247 -691 1299
rect -639 1247 -626 1299
rect -574 1247 -562 1299
rect -510 1247 -498 1299
rect -446 1247 -434 1299
rect -382 1247 -370 1299
rect -318 1247 -306 1299
rect -254 1247 -242 1299
rect -190 1247 -178 1299
rect -126 1247 -114 1299
rect -62 1247 -50 1299
rect 2 1247 14 1299
rect 66 1247 78 1299
rect 130 1247 142 1299
rect 194 1247 206 1299
rect 258 1247 270 1299
rect 322 1247 334 1299
rect 386 1247 398 1299
rect 450 1247 462 1299
rect 514 1247 526 1299
rect 578 1247 590 1299
rect 642 1247 654 1299
rect 706 1247 712 1299
rect 5398 1258 5407 1314
rect 5463 1258 5487 1314
rect 5543 1258 5552 1314
rect 22727 1293 22769 1325
tri 24297 1323 24299 1325 se
rect 24299 1323 24347 1325
tri 24347 1323 24385 1361 nw
tri 24289 1315 24297 1323 se
rect 24297 1315 24333 1323
tri 24288 1314 24289 1315 se
rect 24289 1314 24333 1315
tri 24283 1309 24288 1314 se
rect 24288 1309 24333 1314
tri 24333 1309 24347 1323 nw
tri 24271 1297 24283 1309 se
rect 24283 1297 24321 1309
tri 24321 1297 24333 1309 nw
tri 24267 1293 24271 1297 se
rect 24271 1293 24315 1297
tri 24265 1291 24267 1293 se
rect 24267 1291 24315 1293
tri 24315 1291 24321 1297 nw
tri 24247 1273 24265 1291 se
rect 24265 1273 24297 1291
tri 24297 1273 24315 1291 nw
tri 24232 1258 24247 1273 se
rect 24247 1258 24264 1273
rect -892 1227 712 1247
rect -892 1175 -886 1227
rect -834 1175 -821 1227
rect -769 1175 -756 1227
rect -704 1175 -691 1227
rect -639 1175 -626 1227
rect -574 1175 -562 1227
rect -510 1175 -498 1227
rect -446 1175 -434 1227
rect -382 1175 -370 1227
rect -318 1175 -306 1227
rect -254 1175 -242 1227
rect -190 1175 -178 1227
rect -126 1175 -114 1227
rect -62 1175 -50 1227
rect 2 1175 14 1227
rect 66 1175 78 1227
rect 130 1175 142 1227
rect 194 1175 206 1227
rect 258 1175 270 1227
rect 322 1175 334 1227
rect 386 1175 398 1227
rect 450 1175 462 1227
rect 514 1175 526 1227
rect 578 1175 590 1227
rect 642 1175 654 1227
rect 706 1175 712 1227
tri 24214 1240 24232 1258 se
rect 24232 1240 24264 1258
tri 24264 1240 24297 1273 nw
tri 24476 1253 24490 1267 se
rect 24490 1253 24522 2998
rect 24614 2718 24801 2724
rect 24666 2666 24801 2718
rect 24614 2653 24801 2666
rect 24666 2601 24801 2653
rect 24614 2595 24801 2601
tri 24715 2561 24749 2595 ne
rect 24578 1447 24584 1499
rect 24636 1447 24649 1499
rect 24701 1447 24707 1499
tri 24621 1413 24655 1447 ne
tri 24465 1242 24476 1253 se
rect 24476 1242 24511 1253
tri 24511 1242 24522 1253 nw
tri 24463 1240 24465 1242 se
rect 24465 1240 24509 1242
tri 24509 1240 24511 1242 nw
rect 24214 1239 24263 1240
tri 24263 1239 24264 1240 nw
tri 24462 1239 24463 1240 se
rect 24463 1239 24508 1240
tri 24508 1239 24509 1240 nw
rect 24214 1226 24250 1239
tri 24250 1226 24263 1239 nw
tri 24449 1226 24462 1239 se
rect 24462 1226 24495 1239
tri 24495 1226 24508 1239 nw
rect -892 1155 712 1175
rect 5963 1170 5972 1226
rect 6028 1170 6052 1226
rect 6108 1170 6117 1226
rect -892 1103 -886 1155
rect -834 1103 -821 1155
rect -769 1103 -756 1155
rect -704 1103 -691 1155
rect -639 1103 -626 1155
rect -574 1103 -562 1155
rect -510 1103 -498 1155
rect -446 1103 -434 1155
rect -382 1103 -370 1155
rect -318 1103 -306 1155
rect -254 1103 -242 1155
rect -190 1103 -178 1155
rect -126 1103 -114 1155
rect -62 1103 -50 1155
rect 2 1103 14 1155
rect 66 1103 78 1155
rect 130 1103 142 1155
rect 194 1103 206 1155
rect 258 1103 270 1155
rect 322 1103 334 1155
rect 386 1103 398 1155
rect 450 1103 462 1155
rect 514 1103 526 1155
rect 578 1103 590 1155
rect 642 1103 654 1155
rect 706 1103 712 1155
rect 18784 1126 18964 1132
rect -892 1083 712 1103
rect 16971 1099 17027 1108
rect -892 1031 -886 1083
rect -834 1031 -821 1083
rect -769 1031 -756 1083
rect -704 1031 -691 1083
rect -639 1031 -626 1083
rect -574 1031 -562 1083
rect -510 1031 -498 1083
rect -446 1031 -434 1083
rect -382 1031 -370 1083
rect -318 1031 -306 1083
rect -254 1031 -242 1083
rect -190 1031 -178 1083
rect -126 1031 -114 1083
rect -62 1031 -50 1083
rect 2 1031 14 1083
rect 66 1031 78 1083
rect 130 1031 142 1083
rect 194 1031 206 1083
rect 258 1031 270 1083
rect 322 1031 334 1083
rect 386 1031 398 1083
rect 450 1031 462 1083
rect 514 1031 526 1083
rect 578 1031 590 1083
rect 642 1031 654 1083
rect 706 1031 712 1083
rect -892 1011 712 1031
rect -892 959 -886 1011
rect -834 959 -821 1011
rect -769 959 -756 1011
rect -704 959 -691 1011
rect -639 959 -626 1011
rect -574 959 -562 1011
rect -510 959 -498 1011
rect -446 959 -434 1011
rect -382 959 -370 1011
rect -318 959 -306 1011
rect -254 959 -242 1011
rect -190 959 -178 1011
rect -126 959 -114 1011
rect -62 959 -50 1011
rect 2 959 14 1011
rect 66 959 78 1011
rect 130 959 142 1011
rect 194 959 206 1011
rect 258 959 270 1011
rect 322 959 334 1011
rect 386 959 398 1011
rect 450 959 462 1011
rect 514 959 526 1011
rect 578 959 590 1011
rect 642 959 654 1011
rect 706 959 712 1011
rect -892 939 712 959
rect -892 887 -886 939
rect -834 887 -821 939
rect -769 887 -756 939
rect -704 887 -691 939
rect -639 887 -626 939
rect -574 887 -562 939
rect -510 887 -498 939
rect -446 887 -434 939
rect -382 887 -370 939
rect -318 887 -306 939
rect -254 887 -242 939
rect -190 887 -178 939
rect -126 887 -114 939
rect -62 887 -50 939
rect 2 887 14 939
rect 66 887 78 939
rect 130 887 142 939
rect 194 887 206 939
rect 258 887 270 939
rect 322 887 334 939
rect 386 887 398 939
rect 450 887 462 939
rect 514 887 526 939
rect 578 887 590 939
rect 642 887 654 939
rect 706 887 712 939
rect 7857 1074 7993 1083
rect 18985 1066 19010 1122
rect 19066 1066 19075 1122
rect 17547 1054 17642 1055
rect 16971 1019 17027 1043
rect 16971 954 17027 963
rect 17491 1045 17642 1054
rect 17547 989 17642 1045
rect 17491 965 17642 989
rect 7857 929 7993 938
rect 17547 909 17642 965
rect 18964 996 19075 1066
tri 23943 1036 23948 1041 se
rect 23948 1036 23954 1041
rect 18784 940 18848 946
rect 18904 940 18929 946
rect 18985 940 19010 996
rect 19066 940 19075 996
tri 23359 989 23406 1036 se
rect 23406 989 23954 1036
rect 24006 989 24019 1041
rect 24071 989 24077 1041
tri 23336 966 23359 989 se
rect 23359 966 23406 989
tri 23406 966 23429 989 nw
tri 24203 966 24214 977 se
rect 24214 966 24242 1226
tri 24242 1218 24250 1226 nw
tri 24441 1218 24449 1226 se
rect 24449 1218 24487 1226
tri 24487 1218 24495 1226 nw
tri 24433 1210 24441 1218 se
rect 24441 1210 24465 1218
tri 23331 961 23336 966 se
rect 23336 961 23401 966
tri 23401 961 23406 966 nw
tri 24198 961 24203 966 se
rect 24203 961 24242 966
tri 24417 961 24433 977 se
rect 24433 961 24465 1210
tri 24465 1196 24487 1218 nw
tri 24639 961 24655 977 se
rect 24655 961 24707 1447
rect 24749 1120 24801 2595
rect 25325 1730 25377 5044
rect 25416 5156 25468 5184
rect 25416 1813 25468 5104
tri 25416 1774 25455 1813 ne
rect 25455 1774 25468 1813
tri 25468 1774 25520 1826 sw
tri 25455 1765 25464 1774 ne
rect 25464 1765 25520 1774
tri 25520 1765 25529 1774 sw
tri 25377 1730 25412 1765 sw
tri 25464 1761 25468 1765 ne
rect 25468 1761 25529 1765
tri 25468 1730 25499 1761 ne
rect 25499 1730 25529 1761
tri 25529 1730 25564 1765 sw
rect 25325 1722 25412 1730
tri 25325 1635 25412 1722 ne
tri 25412 1709 25433 1730 sw
tri 25499 1709 25520 1730 ne
rect 25520 1709 25564 1730
tri 25564 1709 25585 1730 sw
rect 25412 1635 25433 1709
tri 25433 1635 25507 1709 sw
tri 25520 1644 25585 1709 ne
tri 25585 1644 25650 1709 sw
tri 25585 1635 25594 1644 ne
rect 25594 1635 25650 1644
tri 25650 1635 25659 1644 sw
tri 25412 1600 25447 1635 ne
rect 25447 1600 25507 1635
tri 25507 1600 25542 1635 sw
tri 25594 1600 25629 1635 ne
rect 25629 1600 25659 1635
tri 25659 1600 25694 1635 sw
tri 25447 1576 25471 1600 ne
rect 25471 1576 25542 1600
tri 25542 1576 25566 1600 sw
tri 25629 1579 25650 1600 ne
rect 25650 1579 25694 1600
tri 25694 1579 25715 1600 sw
tri 25650 1576 25653 1579 ne
rect 25653 1576 25715 1579
tri 25715 1576 25718 1579 sw
tri 25471 1540 25507 1576 ne
rect 25507 1540 25566 1576
tri 25566 1540 25602 1576 sw
tri 25653 1540 25689 1576 ne
rect 25689 1540 25718 1576
tri 25718 1540 25754 1576 sw
tri 25507 1445 25602 1540 ne
tri 25602 1514 25628 1540 sw
tri 25689 1514 25715 1540 ne
rect 25715 1514 25754 1540
tri 25754 1514 25780 1540 sw
rect 25602 1445 25628 1514
tri 25628 1445 25697 1514 sw
tri 25715 1501 25728 1514 ne
tri 25602 1402 25645 1445 ne
rect 25095 1239 25101 1291
rect 25153 1239 25165 1291
rect 25217 1239 25223 1291
tri 25100 1205 25134 1239 ne
tri 24801 1120 24835 1154 sw
rect 24749 1068 24755 1120
rect 24807 1068 24819 1120
rect 24871 1068 24877 1120
tri 24707 961 24723 977 sw
tri 23313 943 23331 961 se
rect 23331 943 23383 961
tri 23383 943 23401 961 nw
tri 24180 943 24198 961 se
rect 24198 943 24242 961
tri 24399 943 24417 961 se
rect 24417 943 24465 961
tri 24621 943 24639 961 se
rect 24639 943 24723 961
tri 24723 943 24741 961 sw
tri 23310 940 23313 943 se
rect 23313 940 23378 943
rect 17491 901 17642 909
tri 23308 938 23310 940 se
rect 23310 938 23378 940
tri 23378 938 23383 943 nw
rect 17491 900 17547 901
rect -892 867 712 887
rect -892 815 -886 867
rect -834 815 -821 867
rect -769 815 -756 867
rect -704 815 -691 867
rect -639 815 -626 867
rect -574 815 -562 867
rect -510 815 -498 867
rect -446 815 -434 867
rect -382 815 -370 867
rect -318 815 -306 867
rect -254 815 -242 867
rect -190 815 -178 867
rect -126 815 -114 867
rect -62 815 -50 867
rect 2 815 14 867
rect 66 815 78 867
rect 130 815 142 867
rect 194 815 206 867
rect 258 815 270 867
rect 322 815 334 867
rect 386 815 398 867
rect 450 815 462 867
rect 514 815 526 867
rect 578 815 590 867
rect 642 815 654 867
rect 706 815 712 867
rect -892 813 712 815
tri 23294 563 23308 577 se
rect 23308 563 23358 938
tri 23358 918 23378 938 nw
rect 24051 891 24057 943
rect 24109 891 24121 943
rect 24173 891 24242 943
rect 24337 891 24343 943
rect 24395 891 24407 943
rect 24459 891 24465 943
rect 24618 891 24624 943
rect 24676 891 24688 943
rect 24740 891 24746 943
rect 24925 909 24931 961
rect 24983 909 24995 961
rect 25047 909 25053 961
tri 25112 911 25134 933 se
rect 25134 911 25186 1239
tri 25186 1205 25220 1239 nw
tri 25186 911 25208 933 sw
rect 25645 911 25697 1445
rect 25728 1361 25780 1514
rect 25728 1297 25780 1309
rect 25728 1239 25780 1245
tri 25110 909 25112 911 se
rect 25112 909 25208 911
rect 24925 899 25001 909
tri 25001 899 25011 909 nw
tri 25100 899 25110 909 se
rect 25110 899 25208 909
tri 25208 899 25220 911 sw
tri 24891 741 24925 775 se
rect 24925 741 24977 899
tri 24977 875 25001 899 nw
rect 25095 847 25101 899
rect 25153 847 25165 899
rect 25217 847 25223 899
rect 25645 847 25697 859
rect 25645 787 25697 795
rect 24827 689 24833 741
rect 24885 718 24897 741
rect 24949 689 24977 741
tri 24841 659 24871 689 ne
rect 24871 662 24875 689
rect 24871 659 24931 662
rect 24501 650 24557 659
tri 24871 655 24875 659 ne
tri 23358 563 23375 580 sw
rect 24501 570 24557 594
rect 24875 638 24931 659
tri 24931 655 24965 689 nw
rect 24875 573 24931 582
tri 23277 546 23294 563 se
rect 23294 546 23375 563
tri 23375 546 23392 563 sw
rect 23277 494 23283 546
rect 23335 494 23347 546
rect 23399 494 23405 546
rect 24553 511 24557 514
rect 24501 505 24557 511
tri 23207 367 23241 401 se
tri 23224 298 23241 315 ne
rect -730 219 -678 225
rect -253 177 -247 229
rect -195 177 -183 229
rect -131 227 -125 229
rect -131 193 1787 227
rect -131 177 -125 193
rect -730 155 -678 167
rect -730 97 -678 103
rect 1753 48 1787 193
rect 15980 125 17587 140
rect 19407 129 19413 181
rect 19465 129 19477 181
rect 19529 129 19535 181
rect 19407 125 19441 129
rect 11284 106 19441 125
rect 11284 91 16014 106
rect 17553 91 19441 106
rect 11284 56 11318 91
rect 17322 61 17331 78
rect 1753 14 6284 48
rect 5918 -80 5927 -24
rect 5983 -80 6007 -24
rect 6063 -48 6072 -24
rect 6063 -80 6216 -48
rect 6184 -269 6216 -80
rect 6250 -112 6284 14
rect 8201 22 11318 56
rect 11367 29 17331 61
rect 8201 -112 8235 22
rect 11367 -11 11399 29
rect 17322 22 17331 29
rect 17387 22 17411 78
rect 17467 22 17476 78
rect 6250 -146 8235 -112
rect 8287 -43 11399 -11
rect 8287 -269 8319 -43
rect 13231 -65 13237 -13
rect 13423 -65 13438 -13
rect 13557 -65 13558 -13
rect 13624 -65 13639 -13
rect 13757 -65 13764 -13
rect 13823 -65 13829 -13
rect 13231 -69 13248 -65
rect 13304 -69 13352 -65
rect 13408 -69 13455 -65
rect 13511 -69 13558 -65
rect 13614 -69 13661 -65
rect 13717 -69 13764 -65
rect 13820 -69 13829 -65
rect 13231 -113 13829 -69
rect 13231 -117 13248 -113
rect 13304 -117 13352 -113
rect 13408 -117 13455 -113
rect 13511 -117 13558 -113
rect 13614 -117 13661 -113
rect 13717 -117 13764 -113
rect 13820 -117 13829 -113
rect 13231 -169 13237 -117
rect 13423 -169 13438 -117
rect 13557 -169 13558 -117
rect 13624 -169 13639 -117
rect 13757 -169 13764 -117
rect 13823 -169 13829 -117
rect 6184 -301 8319 -269
rect 11939 -1733 11976 -1708
rect 24501 -1713 24557 -1704
rect 24501 -1793 24557 -1769
tri 24486 -1814 24501 -1799 se
tri 24356 -1858 24400 -1814 se
rect 24400 -1849 24501 -1814
rect 24400 -1858 24557 -1849
tri 24355 -1859 24356 -1858 se
rect 24356 -1859 24404 -1858
rect 23359 -2001 23415 -1996
rect 24355 -2001 24404 -1859
tri 24404 -1882 24428 -1858 nw
rect 23358 -2005 24404 -2001
rect 23358 -2057 23359 -2005
rect 23415 -2056 24404 -2005
rect 23415 -2057 24398 -2056
rect 23359 -2085 23415 -2061
rect 23359 -2150 23415 -2141
rect 666 -4288 722 -4279
rect 666 -4345 722 -4344
rect 635 -4361 765 -4345
rect 635 -4413 641 -4361
rect 693 -4368 707 -4361
rect 759 -4413 765 -4361
rect 635 -4424 666 -4413
rect 722 -4424 765 -4413
rect 635 -4429 765 -4424
rect 666 -4433 722 -4429
<< via2 >>
rect 8103 7899 8159 7955
rect 8193 7899 8249 7955
rect 8283 7899 8339 7955
rect 8372 7899 8428 7955
rect 8461 7899 8517 7955
rect 8103 7819 8159 7875
rect 8193 7819 8249 7875
rect 8283 7819 8339 7875
rect 8372 7819 8428 7875
rect 8461 7819 8517 7875
rect 6575 7553 6711 7769
rect 8103 7739 8159 7795
rect 8193 7739 8249 7795
rect 8283 7739 8339 7795
rect 8372 7739 8428 7795
rect 8461 7739 8517 7795
rect 12750 7899 12806 7955
rect 12840 7899 12896 7955
rect 12930 7899 12986 7955
rect 13019 7899 13075 7955
rect 13108 7899 13164 7955
rect 12750 7819 12806 7875
rect 12840 7819 12896 7875
rect 12930 7819 12986 7875
rect 13019 7819 13075 7875
rect 13108 7819 13164 7875
rect 12750 7739 12806 7795
rect 12840 7739 12896 7795
rect 12930 7739 12986 7795
rect 13019 7739 13075 7795
rect 13108 7739 13164 7795
rect 14279 7899 14335 7955
rect 14367 7899 14423 7955
rect 14455 7899 14511 7955
rect 14543 7899 14599 7955
rect 14630 7899 14686 7955
rect 14279 7819 14335 7875
rect 14367 7819 14423 7875
rect 14455 7819 14511 7875
rect 14543 7819 14599 7875
rect 14630 7819 14686 7875
rect 14279 7739 14335 7795
rect 14367 7739 14423 7795
rect 14455 7739 14511 7795
rect 14543 7739 14599 7795
rect 14630 7739 14686 7795
rect 15846 7839 15982 8055
rect 8102 5778 8158 5834
rect 8192 5778 8248 5834
rect 8282 5778 8338 5834
rect 8371 5778 8427 5834
rect 8460 5778 8516 5834
rect 14275 5778 14331 5834
rect 14365 5778 14421 5834
rect 14455 5778 14511 5834
rect 14544 5778 14600 5834
rect 14633 5778 14689 5834
rect 8102 5698 8158 5754
rect 8192 5698 8248 5754
rect 8282 5698 8338 5754
rect 8371 5698 8427 5754
rect 8460 5698 8516 5754
rect 14275 5698 14331 5754
rect 14365 5698 14421 5754
rect 14455 5698 14511 5754
rect 14544 5698 14600 5754
rect 14633 5698 14689 5754
rect 15841 5672 15897 5728
rect 15931 5672 15987 5728
rect 17068 5681 17124 5737
rect 17151 5681 17207 5737
rect 17234 5681 17290 5737
rect 12750 5575 12806 5631
rect 12840 5575 12896 5631
rect 12930 5575 12986 5631
rect 13019 5575 13075 5631
rect 13108 5575 13164 5631
rect 15841 5547 15897 5603
rect 15931 5547 15987 5603
rect 17068 5539 17124 5595
rect 17151 5539 17207 5595
rect 17234 5539 17290 5595
rect 11090 5420 11146 5476
rect 11174 5420 11230 5476
rect 11258 5420 11314 5476
rect 11342 5420 11398 5476
rect 13761 5420 13817 5476
rect 13845 5420 13901 5476
rect 13929 5420 13985 5476
rect 14013 5420 14069 5476
rect 12908 4014 12964 4070
rect 5401 3901 5457 3957
rect 5481 3901 5537 3957
rect 12908 3930 12964 3986
rect 16877 3703 16933 3759
rect 16957 3703 17013 3759
rect 17451 3711 17507 3767
rect 17531 3711 17587 3767
rect 12084 3211 12140 3267
rect 12908 3211 12964 3267
rect 10285 3197 10341 3198
rect 10367 3197 10423 3198
rect 10449 3197 10505 3198
rect 10530 3197 10586 3198
rect 10611 3197 10667 3198
rect 10692 3197 10748 3198
rect 10285 3145 10286 3197
rect 10286 3145 10338 3197
rect 10338 3145 10341 3197
rect 10367 3145 10407 3197
rect 10407 3145 10423 3197
rect 10449 3145 10475 3197
rect 10475 3145 10491 3197
rect 10491 3145 10505 3197
rect 10530 3145 10543 3197
rect 10543 3145 10559 3197
rect 10559 3145 10586 3197
rect 10611 3145 10627 3197
rect 10627 3145 10667 3197
rect 10692 3145 10695 3197
rect 10695 3145 10747 3197
rect 10747 3145 10748 3197
rect 10285 3142 10341 3145
rect 10367 3142 10423 3145
rect 10449 3142 10505 3145
rect 10530 3142 10586 3145
rect 10611 3142 10667 3145
rect 10692 3142 10748 3145
rect 12084 3131 12140 3187
rect 12908 3131 12964 3187
rect 10285 3061 10286 3096
rect 10286 3061 10338 3096
rect 10338 3061 10341 3096
rect 10367 3061 10407 3096
rect 10407 3061 10423 3096
rect 10449 3061 10475 3096
rect 10475 3061 10491 3096
rect 10491 3061 10505 3096
rect 10530 3061 10543 3096
rect 10543 3061 10559 3096
rect 10559 3061 10586 3096
rect 10611 3061 10627 3096
rect 10627 3061 10667 3096
rect 10692 3061 10695 3096
rect 10695 3061 10747 3096
rect 10747 3061 10748 3096
rect 10285 3040 10341 3061
rect 10367 3040 10423 3061
rect 10449 3040 10505 3061
rect 10530 3040 10586 3061
rect 10611 3040 10667 3061
rect 10692 3040 10748 3061
rect 17365 2689 17421 2745
rect 17745 2691 17801 2747
rect 17365 2609 17421 2665
rect 17745 2611 17801 2667
rect 20743 2405 20799 2417
rect 20825 2405 20881 2417
rect 20907 2405 20963 2417
rect 20989 2405 21045 2417
rect 21071 2405 21127 2417
rect 20743 2361 20794 2405
rect 20794 2361 20799 2405
rect 20825 2361 20861 2405
rect 20861 2361 20876 2405
rect 20876 2361 20881 2405
rect 20907 2361 20928 2405
rect 20928 2361 20943 2405
rect 20943 2361 20963 2405
rect 20989 2361 20995 2405
rect 20995 2361 21010 2405
rect 21010 2361 21045 2405
rect 21071 2361 21076 2405
rect 21076 2361 21127 2405
rect 20743 2331 20799 2337
rect 20825 2331 20881 2337
rect 20907 2331 20963 2337
rect 20989 2331 21045 2337
rect 21071 2331 21127 2337
rect 18848 2270 18894 2319
rect 18894 2270 18904 2319
rect 18936 2270 18968 2319
rect 18968 2270 18990 2319
rect 18990 2270 18992 2319
rect 19024 2270 19042 2319
rect 19042 2270 19064 2319
rect 19064 2270 19080 2319
rect 19112 2270 19116 2319
rect 19116 2270 19168 2319
rect 18848 2263 18904 2270
rect 18936 2263 18992 2270
rect 19024 2263 19080 2270
rect 19112 2263 19168 2270
rect 18848 2187 18904 2193
rect 18936 2187 18992 2193
rect 19024 2187 19080 2193
rect 19112 2187 19168 2193
rect 18848 2137 18894 2187
rect 18894 2137 18904 2187
rect 18936 2137 18968 2187
rect 18968 2137 18990 2187
rect 18990 2137 18992 2187
rect 19024 2137 19042 2187
rect 19042 2137 19064 2187
rect 19064 2137 19080 2187
rect 19112 2137 19116 2187
rect 19116 2137 19168 2187
rect 20743 2281 20794 2331
rect 20794 2281 20799 2331
rect 20825 2281 20861 2331
rect 20861 2281 20876 2331
rect 20876 2281 20881 2331
rect 20907 2281 20928 2331
rect 20928 2281 20943 2331
rect 20943 2281 20963 2331
rect 20989 2281 20995 2331
rect 20995 2281 21010 2331
rect 21010 2281 21045 2331
rect 21071 2281 21076 2331
rect 21076 2281 21127 2331
rect 20743 2205 20794 2257
rect 20794 2205 20799 2257
rect 20825 2205 20861 2257
rect 20861 2205 20876 2257
rect 20876 2205 20881 2257
rect 20907 2205 20928 2257
rect 20928 2205 20943 2257
rect 20943 2205 20963 2257
rect 20989 2205 20995 2257
rect 20995 2205 21010 2257
rect 21010 2205 21045 2257
rect 21071 2205 21076 2257
rect 21076 2205 21127 2257
rect 20743 2201 20799 2205
rect 20825 2201 20881 2205
rect 20907 2201 20963 2205
rect 20989 2201 21045 2205
rect 21071 2201 21127 2205
rect 20743 2131 20794 2177
rect 20794 2131 20799 2177
rect 20825 2131 20861 2177
rect 20861 2131 20876 2177
rect 20876 2131 20881 2177
rect 20907 2131 20928 2177
rect 20928 2131 20943 2177
rect 20943 2131 20963 2177
rect 20989 2131 20995 2177
rect 20995 2131 21010 2177
rect 21010 2131 21045 2177
rect 21071 2131 21076 2177
rect 21076 2131 21127 2177
rect 20743 2121 20799 2131
rect 20825 2121 20881 2131
rect 20907 2121 20963 2131
rect 20989 2121 21045 2131
rect 21071 2121 21127 2131
rect 20743 2057 20794 2097
rect 20794 2057 20799 2097
rect 20825 2057 20861 2097
rect 20861 2057 20876 2097
rect 20876 2057 20881 2097
rect 20907 2057 20928 2097
rect 20928 2057 20943 2097
rect 20943 2057 20963 2097
rect 20989 2057 20995 2097
rect 20995 2057 21010 2097
rect 21010 2057 21045 2097
rect 21071 2057 21076 2097
rect 21076 2057 21127 2097
rect 20743 2041 20799 2057
rect 20825 2041 20881 2057
rect 20907 2041 20963 2057
rect 20989 2041 21045 2057
rect 21071 2041 21127 2057
rect 10357 1613 10406 1665
rect 10406 1613 10413 1665
rect 10480 1613 10487 1665
rect 10487 1613 10536 1665
rect 10357 1609 10413 1613
rect 10480 1609 10536 1613
rect 10357 1521 10406 1563
rect 10406 1521 10413 1563
rect 10480 1521 10487 1563
rect 10487 1521 10536 1563
rect 10357 1507 10413 1521
rect 10480 1507 10536 1521
rect 12084 1404 12140 1460
rect 12084 1324 12140 1380
rect 5407 1258 5463 1314
rect 5487 1258 5543 1314
rect 5972 1170 6028 1226
rect 6052 1170 6108 1226
rect 7857 938 7993 1074
rect 16971 1043 17027 1099
rect 18848 1066 18904 1122
rect 18929 1066 18964 1122
rect 18964 1066 18985 1122
rect 19010 1066 19066 1122
rect 16971 963 17027 1019
rect 17491 989 17547 1045
rect 17491 909 17547 965
rect 18848 946 18904 996
rect 18929 946 18964 996
rect 18964 946 18985 996
rect 18848 940 18904 946
rect 18929 940 18985 946
rect 19010 940 19066 996
rect 24875 689 24885 718
rect 24885 689 24897 718
rect 24897 689 24931 718
rect 24875 662 24931 689
rect 24501 649 24557 650
rect 24501 597 24553 649
rect 24553 597 24557 649
rect 24501 594 24557 597
rect 24875 582 24931 638
rect 24501 563 24557 570
rect 24501 514 24553 563
rect 24553 514 24557 563
rect 5927 -80 5983 -24
rect 6007 -80 6063 -24
rect 17331 22 17387 78
rect 17411 22 17467 78
rect 13248 -65 13289 -13
rect 13289 -65 13304 -13
rect 13352 -65 13356 -13
rect 13356 -65 13371 -13
rect 13371 -65 13408 -13
rect 13455 -65 13490 -13
rect 13490 -65 13505 -13
rect 13505 -65 13511 -13
rect 13558 -65 13572 -13
rect 13572 -65 13614 -13
rect 13661 -65 13691 -13
rect 13691 -65 13705 -13
rect 13705 -65 13717 -13
rect 13764 -65 13771 -13
rect 13771 -65 13820 -13
rect 13248 -69 13304 -65
rect 13352 -69 13408 -65
rect 13455 -69 13511 -65
rect 13558 -69 13614 -65
rect 13661 -69 13717 -65
rect 13764 -69 13820 -65
rect 13248 -117 13304 -113
rect 13352 -117 13408 -113
rect 13455 -117 13511 -113
rect 13558 -117 13614 -113
rect 13661 -117 13717 -113
rect 13764 -117 13820 -113
rect 13248 -169 13289 -117
rect 13289 -169 13304 -117
rect 13352 -169 13356 -117
rect 13356 -169 13371 -117
rect 13371 -169 13408 -117
rect 13455 -169 13490 -117
rect 13490 -169 13505 -117
rect 13505 -169 13511 -117
rect 13558 -169 13572 -117
rect 13572 -169 13614 -117
rect 13661 -169 13691 -117
rect 13691 -169 13705 -117
rect 13705 -169 13717 -117
rect 13764 -169 13771 -117
rect 13771 -169 13820 -117
rect 24501 -1769 24557 -1713
rect 24501 -1849 24557 -1793
rect 23359 -2061 23415 -2005
rect 23359 -2141 23415 -2085
rect 666 -4344 722 -4288
rect 666 -4413 693 -4368
rect 693 -4413 707 -4368
rect 707 -4413 722 -4368
rect 666 -4424 722 -4413
<< metal3 >>
rect 15841 8055 15987 8060
rect 8098 7955 8522 7960
rect 8098 7899 8103 7955
rect 8159 7899 8193 7955
rect 8249 7899 8283 7955
rect 8339 7899 8372 7955
rect 8428 7899 8461 7955
rect 8517 7899 8522 7955
rect 8098 7875 8522 7899
rect 8098 7819 8103 7875
rect 8159 7819 8193 7875
rect 8249 7819 8283 7875
rect 8339 7819 8372 7875
rect 8428 7819 8461 7875
rect 8517 7819 8522 7875
rect 8098 7795 8522 7819
rect 8098 7774 8103 7795
rect 6570 7769 6716 7774
rect 6570 7553 6575 7769
rect 6711 7553 6716 7769
rect 6570 5384 6716 7553
rect 8097 7739 8103 7774
rect 8159 7739 8193 7795
rect 8249 7739 8283 7795
rect 8339 7739 8372 7795
rect 8428 7739 8461 7795
rect 8517 7739 8522 7795
rect 8097 5834 8522 7739
rect 8097 5778 8102 5834
rect 8158 5778 8192 5834
rect 8248 5778 8282 5834
rect 8338 5778 8371 5834
rect 8427 5778 8460 5834
rect 8516 5778 8522 5834
rect 8097 5754 8522 5778
rect 8097 5698 8102 5754
rect 8158 5698 8192 5754
rect 8248 5698 8282 5754
rect 8338 5698 8371 5754
rect 8427 5698 8460 5754
rect 8516 5703 8522 5754
rect 12745 7955 13169 7960
rect 12745 7899 12750 7955
rect 12806 7899 12840 7955
rect 12896 7899 12930 7955
rect 12986 7899 13019 7955
rect 13075 7899 13108 7955
rect 13164 7899 13169 7955
rect 12745 7875 13169 7899
rect 12745 7819 12750 7875
rect 12806 7819 12840 7875
rect 12896 7819 12930 7875
rect 12986 7819 13019 7875
rect 13075 7819 13108 7875
rect 13164 7819 13169 7875
rect 12745 7795 13169 7819
rect 12745 7739 12750 7795
rect 12806 7739 12840 7795
rect 12896 7739 12930 7795
rect 12986 7739 13019 7795
rect 13075 7739 13108 7795
rect 13164 7739 13169 7795
rect 14274 7955 14691 7960
rect 14274 7899 14279 7955
rect 14335 7899 14367 7955
rect 14423 7899 14455 7955
rect 14511 7899 14543 7955
rect 14599 7899 14630 7955
rect 14686 7899 14691 7955
rect 14274 7875 14691 7899
rect 14274 7819 14279 7875
rect 14335 7819 14367 7875
rect 14423 7819 14455 7875
rect 14511 7819 14543 7875
rect 14599 7819 14630 7875
rect 14686 7819 14691 7875
rect 14274 7795 14691 7819
rect 14274 7774 14279 7795
rect 8516 5698 8521 5703
rect 8097 5693 8521 5698
rect 12745 5631 13169 7739
rect 14270 7739 14279 7774
rect 14335 7739 14367 7795
rect 14423 7739 14455 7795
rect 14511 7739 14543 7795
rect 14599 7739 14630 7795
rect 14686 7774 14691 7795
rect 15841 7839 15846 8055
rect 15982 7839 15987 8055
rect 14686 7739 14695 7774
rect 14270 5834 14695 7739
rect 14270 5778 14275 5834
rect 14331 5778 14365 5834
rect 14421 5778 14455 5834
rect 14511 5778 14544 5834
rect 14600 5778 14633 5834
rect 14689 5778 14695 5834
rect 14270 5754 14695 5778
rect 14270 5698 14275 5754
rect 14331 5698 14365 5754
rect 14421 5698 14455 5754
rect 14511 5698 14544 5754
rect 14600 5698 14633 5754
rect 14689 5703 14695 5754
rect 15841 5737 15987 7839
rect 17059 5737 17299 5742
rect 15836 5728 15992 5737
rect 14689 5698 14694 5703
rect 14270 5693 14694 5698
rect 12745 5575 12750 5631
rect 12806 5575 12840 5631
rect 12896 5575 12930 5631
rect 12986 5575 13019 5631
rect 13075 5575 13108 5631
rect 13164 5575 13169 5631
rect 12745 5539 13169 5575
rect 15836 5672 15841 5728
rect 15897 5672 15931 5728
rect 15987 5672 15992 5728
rect 15836 5603 15992 5672
rect 15836 5547 15841 5603
rect 15897 5547 15931 5603
rect 15987 5547 15992 5603
rect 15836 5538 15992 5547
rect 17059 5681 17068 5737
rect 17124 5681 17151 5737
rect 17207 5681 17234 5737
rect 17290 5681 17299 5737
rect 17059 5595 17299 5681
rect 17059 5539 17068 5595
rect 17124 5539 17151 5595
rect 17207 5539 17234 5595
rect 17290 5539 17299 5595
rect 11085 5476 11403 5512
rect 11085 5420 11090 5476
rect 11146 5420 11174 5476
rect 11230 5420 11258 5476
rect 11314 5420 11342 5476
rect 11398 5420 11403 5476
tri 6716 5384 6731 5399 sw
rect 11085 5384 11403 5420
rect 13756 5476 14074 5512
rect 13756 5420 13761 5476
rect 13817 5420 13845 5476
rect 13901 5420 13929 5476
rect 13985 5420 14013 5476
rect 14069 5420 14074 5476
rect 13756 5384 14074 5420
rect 6570 5214 6731 5384
tri 6731 5214 6901 5384 sw
rect 6570 5205 6901 5214
tri 6570 5096 6679 5205 ne
rect 6679 5096 6901 5205
rect 17059 5096 17299 5539
rect 20734 5504 21132 5516
rect 20734 5440 20740 5504
rect 20804 5440 20820 5504
rect 20884 5440 20900 5504
rect 20964 5440 20980 5504
rect 21044 5440 21060 5504
rect 21124 5440 21132 5504
rect 20734 5418 21132 5440
rect 20734 5354 20740 5418
rect 20804 5354 20820 5418
rect 20884 5354 20900 5418
rect 20964 5354 20980 5418
rect 21044 5354 21060 5418
rect 21124 5354 21132 5418
rect 20734 5332 21132 5354
rect 20734 5268 20740 5332
rect 20804 5268 20820 5332
rect 20884 5268 20900 5332
rect 20964 5268 20980 5332
rect 21044 5268 21060 5332
rect 21124 5268 21132 5332
rect 20734 5246 21132 5268
rect 20734 5182 20740 5246
rect 20804 5182 20820 5246
rect 20884 5182 20900 5246
rect 20964 5182 20980 5246
rect 21044 5182 21060 5246
rect 21124 5182 21132 5246
rect 20734 5160 21132 5182
rect 20734 5096 20740 5160
rect 20804 5096 20820 5160
rect 20884 5096 20900 5160
rect 20964 5096 20980 5160
rect 21044 5096 21060 5160
rect 21124 5096 21132 5160
tri 6679 5080 6695 5096 ne
rect 6695 5080 6901 5096
rect 20734 5074 21132 5096
rect 20734 5010 20740 5074
rect 20804 5010 20820 5074
rect 20884 5010 20900 5074
rect 20964 5010 20980 5074
rect 21044 5010 21060 5074
rect 21124 5010 21132 5074
rect 20734 4988 21132 5010
rect 20734 4924 20740 4988
rect 20804 4924 20820 4988
rect 20884 4924 20900 4988
rect 20964 4924 20980 4988
rect 21044 4924 21060 4988
rect 21124 4924 21132 4988
rect 20734 4902 21132 4924
rect 20734 4838 20740 4902
rect 20804 4838 20820 4902
rect 20884 4838 20900 4902
rect 20964 4838 20980 4902
rect 21044 4838 21060 4902
rect 21124 4838 21132 4902
rect 20734 4815 21132 4838
rect 20734 4751 20740 4815
rect 20804 4751 20820 4815
rect 20884 4751 20900 4815
rect 20964 4751 20980 4815
rect 21044 4751 21060 4815
rect 21124 4751 21132 4815
rect 20734 4728 21132 4751
rect 20734 4664 20740 4728
rect 20804 4664 20820 4728
rect 20884 4664 20900 4728
rect 20964 4664 20980 4728
rect 21044 4664 21060 4728
rect 21124 4664 21132 4728
rect 11079 4389 11408 4456
rect 13752 4424 14081 4568
rect 12897 4070 12975 4079
rect 12897 4014 12908 4070
rect 12964 4014 12975 4070
rect 12897 3986 12975 4014
rect 5396 3957 5542 3962
rect 5396 3901 5401 3957
rect 5457 3901 5481 3957
rect 5537 3901 5542 3957
rect 12897 3930 12908 3986
rect 12964 3930 12975 3986
rect 12897 3921 12975 3930
rect 5396 3896 5542 3901
tri 5407 1324 5444 1361 se
rect 5444 1324 5510 3896
rect 12078 3267 12147 3276
rect 12078 3211 12084 3267
rect 12140 3211 12147 3267
rect 10217 3198 10817 3203
rect 10217 3142 10285 3198
rect 10341 3142 10367 3198
rect 10423 3142 10449 3198
rect 10505 3142 10530 3198
rect 10586 3142 10611 3198
rect 10667 3142 10692 3198
rect 10748 3142 10817 3198
rect 10217 3096 10817 3142
rect 6602 3053 6856 3061
rect 6441 3049 7070 3053
rect 6441 2985 6447 3049
rect 6511 2985 6540 3049
rect 6604 2985 6632 3049
rect 6696 2985 6724 3049
rect 6788 2985 6816 3049
rect 6880 2985 6908 3049
rect 6972 2985 7000 3049
rect 7064 2985 7070 3049
rect 6441 2963 7070 2985
rect 6441 2899 6447 2963
rect 6511 2899 6540 2963
rect 6604 2899 6632 2963
rect 6696 2899 6724 2963
rect 6788 2899 6816 2963
rect 6880 2899 6908 2963
rect 6972 2899 7000 2963
rect 7064 2899 7070 2963
rect 6441 2877 7070 2899
rect 6441 2813 6447 2877
rect 6511 2813 6540 2877
rect 6604 2813 6632 2877
rect 6696 2813 6724 2877
rect 6788 2813 6816 2877
rect 6880 2813 6908 2877
rect 6972 2813 7000 2877
rect 7064 2813 7070 2877
rect 6441 2791 7070 2813
rect 6441 2727 6447 2791
rect 6511 2727 6540 2791
rect 6604 2727 6632 2791
rect 6696 2727 6724 2791
rect 6788 2727 6816 2791
rect 6880 2727 6908 2791
rect 6972 2727 7000 2791
rect 7064 2727 7070 2791
rect 6441 2705 7070 2727
rect 6441 2641 6447 2705
rect 6511 2641 6540 2705
rect 6604 2641 6632 2705
rect 6696 2641 6724 2705
rect 6788 2641 6816 2705
rect 6880 2641 6908 2705
rect 6972 2641 7000 2705
rect 7064 2641 7070 2705
rect 6441 2619 7070 2641
rect 6441 2555 6447 2619
rect 6511 2555 6540 2619
rect 6604 2555 6632 2619
rect 6696 2555 6724 2619
rect 6788 2555 6816 2619
rect 6880 2555 6908 2619
rect 6972 2555 7000 2619
rect 7064 2555 7070 2619
rect 6441 2533 7070 2555
rect 6441 2469 6447 2533
rect 6511 2469 6540 2533
rect 6604 2469 6632 2533
rect 6696 2469 6724 2533
rect 6788 2469 6816 2533
rect 6880 2469 6908 2533
rect 6972 2469 7000 2533
rect 7064 2469 7070 2533
rect 6441 2465 7070 2469
rect 7869 3049 8504 3053
rect 7869 2985 7875 3049
rect 7939 2985 7969 3049
rect 8033 2985 8062 3049
rect 8126 2985 8155 3049
rect 8219 2985 8248 3049
rect 8312 2985 8341 3049
rect 8405 2985 8434 3049
rect 8498 2985 8504 3049
rect 7869 2963 8504 2985
rect 7869 2899 7875 2963
rect 7939 2899 7969 2963
rect 8033 2899 8062 2963
rect 8126 2899 8155 2963
rect 8219 2899 8248 2963
rect 8312 2899 8341 2963
rect 8405 2899 8434 2963
rect 8498 2899 8504 2963
rect 7869 2877 8504 2899
rect 7869 2813 7875 2877
rect 7939 2813 7969 2877
rect 8033 2813 8062 2877
rect 8126 2813 8155 2877
rect 8219 2813 8248 2877
rect 8312 2813 8341 2877
rect 8405 2813 8434 2877
rect 8498 2813 8504 2877
rect 7869 2791 8504 2813
rect 7869 2727 7875 2791
rect 7939 2727 7969 2791
rect 8033 2727 8062 2791
rect 8126 2727 8155 2791
rect 8219 2727 8248 2791
rect 8312 2727 8341 2791
rect 8405 2727 8434 2791
rect 8498 2727 8504 2791
rect 7869 2705 8504 2727
rect 7869 2641 7875 2705
rect 7939 2641 7969 2705
rect 8033 2641 8062 2705
rect 8126 2641 8155 2705
rect 8219 2641 8248 2705
rect 8312 2641 8341 2705
rect 8405 2641 8434 2705
rect 8498 2641 8504 2705
rect 7869 2619 8504 2641
rect 7869 2555 7875 2619
rect 7939 2555 7969 2619
rect 8033 2555 8062 2619
rect 8126 2555 8155 2619
rect 8219 2555 8248 2619
rect 8312 2555 8341 2619
rect 8405 2555 8434 2619
rect 8498 2555 8504 2619
rect 7869 2533 8504 2555
rect 7869 2469 7875 2533
rect 7939 2469 7969 2533
rect 8033 2469 8062 2533
rect 8126 2469 8155 2533
rect 8219 2469 8248 2533
rect 8312 2469 8341 2533
rect 8405 2469 8434 2533
rect 8498 2469 8504 2533
rect 7869 2465 8504 2469
rect 10217 3040 10285 3096
rect 10341 3040 10367 3096
rect 10423 3040 10449 3096
rect 10505 3040 10530 3096
rect 10586 3040 10611 3096
rect 10667 3040 10692 3096
rect 10748 3040 10817 3096
rect 10217 1665 10817 3040
rect 10217 1609 10357 1665
rect 10413 1609 10480 1665
rect 10536 1609 10817 1665
rect 10217 1563 10817 1609
rect 10217 1507 10357 1563
rect 10413 1507 10480 1563
rect 10536 1507 10817 1563
tri 5510 1324 5547 1361 sw
tri 5406 1323 5407 1324 se
rect 5407 1323 5547 1324
tri 5547 1323 5548 1324 sw
tri 5402 1319 5406 1323 se
rect 5406 1319 5548 1323
rect 5402 1314 5548 1319
rect 5402 1258 5407 1314
rect 5463 1258 5487 1314
rect 5543 1258 5548 1314
rect 5402 1253 5548 1258
rect 5967 1226 6113 1231
rect 5967 1170 5972 1226
rect 6028 1170 6052 1226
rect 6108 1170 6113 1226
rect 5967 1165 6113 1170
rect 6004 -19 6070 1165
rect 10217 1083 10817 1507
rect 12078 3187 12147 3211
rect 12078 3131 12084 3187
rect 12140 3131 12147 3187
rect 12078 1460 12147 3131
rect 12901 3267 12970 3921
rect 17446 3767 17592 3772
rect 16872 3759 17018 3764
rect 16872 3703 16877 3759
rect 16933 3703 16957 3759
rect 17013 3703 17018 3759
rect 17446 3711 17451 3767
rect 17507 3711 17531 3767
rect 17587 3711 17592 3767
rect 17446 3706 17592 3711
rect 16872 3698 17018 3703
rect 12901 3211 12908 3267
rect 12964 3211 12970 3267
rect 12901 3187 12970 3211
rect 12901 3131 12908 3187
rect 12964 3131 12970 3187
rect 12901 3126 12970 3131
rect 16060 2200 16314 2796
rect 15879 2098 16508 2102
rect 15879 2034 15885 2098
rect 15949 2034 15978 2098
rect 16042 2034 16070 2098
rect 16134 2034 16162 2098
rect 16226 2034 16254 2098
rect 16318 2034 16346 2098
rect 16410 2034 16438 2098
rect 16502 2034 16508 2098
rect 15879 2012 16508 2034
rect 15879 1948 15885 2012
rect 15949 1948 15978 2012
rect 16042 1948 16070 2012
rect 16134 1948 16162 2012
rect 16226 1948 16254 2012
rect 16318 1948 16346 2012
rect 16410 1948 16438 2012
rect 16502 1948 16508 2012
rect 15879 1926 16508 1948
rect 15879 1862 15885 1926
rect 15949 1862 15978 1926
rect 16042 1862 16070 1926
rect 16134 1862 16162 1926
rect 16226 1862 16254 1926
rect 16318 1862 16346 1926
rect 16410 1862 16438 1926
rect 16502 1862 16508 1926
rect 15879 1840 16508 1862
rect 15879 1776 15885 1840
rect 15949 1776 15978 1840
rect 16042 1776 16070 1840
rect 16134 1776 16162 1840
rect 16226 1776 16254 1840
rect 16318 1776 16346 1840
rect 16410 1776 16438 1840
rect 16502 1776 16508 1840
rect 15879 1754 16508 1776
rect 15879 1690 15885 1754
rect 15949 1690 15978 1754
rect 16042 1690 16070 1754
rect 16134 1690 16162 1754
rect 16226 1690 16254 1754
rect 16318 1690 16346 1754
rect 16410 1690 16438 1754
rect 16502 1690 16508 1754
rect 15879 1668 16508 1690
rect 15879 1604 15885 1668
rect 15949 1604 15978 1668
rect 16042 1604 16070 1668
rect 16134 1604 16162 1668
rect 16226 1604 16254 1668
rect 16318 1604 16346 1668
rect 16410 1604 16438 1668
rect 16502 1604 16508 1668
rect 15879 1582 16508 1604
rect 15879 1518 15885 1582
rect 15949 1518 15978 1582
rect 16042 1518 16070 1582
rect 16134 1518 16162 1582
rect 16226 1518 16254 1582
rect 16318 1518 16346 1582
rect 16410 1518 16438 1582
rect 16502 1518 16508 1582
rect 15879 1514 16508 1518
rect 12078 1404 12084 1460
rect 12140 1404 12147 1460
rect 12078 1380 12147 1404
rect 12078 1324 12084 1380
rect 12140 1324 12147 1380
rect 12078 1319 12147 1324
rect 16957 1104 17018 3698
rect 17360 2745 17426 2756
rect 17360 2689 17365 2745
rect 17421 2689 17426 2745
rect 17360 2665 17426 2689
rect 17360 2609 17365 2665
rect 17421 2609 17426 2665
rect 16957 1099 17032 1104
rect 5922 -24 6070 -19
rect 5922 -80 5927 -24
rect 5983 -80 6007 -24
rect 6063 -80 6070 -24
rect 5922 -85 6070 -80
rect 7852 1074 7998 1079
rect 7852 938 7857 1074
rect 7993 938 7998 1074
rect 16957 1043 16971 1099
rect 17027 1043 17032 1099
rect 16957 1019 17032 1043
rect 16957 963 16971 1019
rect 17027 963 17032 1019
rect 16957 958 17032 963
tri 7639 -409 7852 -196 se
rect 7852 -263 7998 938
tri 17345 83 17360 98 se
rect 17360 83 17426 2609
rect 17486 1050 17547 3706
rect 17740 2747 17806 3592
rect 17740 2691 17745 2747
rect 17801 2691 17806 2747
rect 17740 2667 17806 2691
rect 17740 2611 17745 2667
rect 17801 2611 17806 2667
rect 17740 2604 17806 2611
rect 20734 2417 21132 4664
rect 20734 2361 20743 2417
rect 20799 2361 20825 2417
rect 20881 2361 20907 2417
rect 20963 2361 20989 2417
rect 21045 2361 21071 2417
rect 21127 2361 21132 2417
rect 20734 2337 21132 2361
rect 18843 2319 19173 2324
rect 18843 2263 18848 2319
rect 18904 2263 18936 2319
rect 18992 2263 19024 2319
rect 19080 2263 19112 2319
rect 19168 2263 19173 2319
rect 18843 2193 19173 2263
rect 18843 2137 18848 2193
rect 18904 2137 18936 2193
rect 18992 2137 19024 2193
rect 19080 2137 19112 2193
rect 19168 2137 19173 2193
rect 18843 2132 19173 2137
rect 20734 2281 20743 2337
rect 20799 2281 20825 2337
rect 20881 2281 20907 2337
rect 20963 2281 20989 2337
rect 21045 2281 21071 2337
rect 21127 2281 21132 2337
rect 20734 2257 21132 2281
rect 20734 2201 20743 2257
rect 20799 2201 20825 2257
rect 20881 2201 20907 2257
rect 20963 2201 20989 2257
rect 21045 2201 21071 2257
rect 21127 2201 21132 2257
rect 20734 2177 21132 2201
rect 20734 2121 20743 2177
rect 20799 2121 20825 2177
rect 20881 2121 20907 2177
rect 20963 2121 20989 2177
rect 21045 2121 21071 2177
rect 21127 2121 21132 2177
rect 17675 2098 18660 2102
rect 17675 2034 17681 2098
rect 17745 2034 17764 2098
rect 17828 2034 17847 2098
rect 17911 2034 17930 2098
rect 17994 2034 18013 2098
rect 18077 2034 18096 2098
rect 18160 2034 18179 2098
rect 18243 2034 18262 2098
rect 18326 2034 18344 2098
rect 18408 2034 18426 2098
rect 18490 2034 18508 2098
rect 18572 2034 18590 2098
rect 18654 2034 18660 2098
rect 17675 2012 18660 2034
rect 17675 1948 17681 2012
rect 17745 1948 17764 2012
rect 17828 1948 17847 2012
rect 17911 1948 17930 2012
rect 17994 1948 18013 2012
rect 18077 1948 18096 2012
rect 18160 1948 18179 2012
rect 18243 1948 18262 2012
rect 18326 1948 18344 2012
rect 18408 1948 18426 2012
rect 18490 1948 18508 2012
rect 18572 1948 18590 2012
rect 18654 1948 18660 2012
rect 17675 1926 18660 1948
rect 17675 1862 17681 1926
rect 17745 1862 17764 1926
rect 17828 1862 17847 1926
rect 17911 1862 17930 1926
rect 17994 1862 18013 1926
rect 18077 1862 18096 1926
rect 18160 1862 18179 1926
rect 18243 1862 18262 1926
rect 18326 1862 18344 1926
rect 18408 1862 18426 1926
rect 18490 1862 18508 1926
rect 18572 1862 18590 1926
rect 18654 1862 18660 1926
rect 17675 1840 18660 1862
rect 17675 1776 17681 1840
rect 17745 1776 17764 1840
rect 17828 1776 17847 1840
rect 17911 1776 17930 1840
rect 17994 1776 18013 1840
rect 18077 1776 18096 1840
rect 18160 1776 18179 1840
rect 18243 1776 18262 1840
rect 18326 1776 18344 1840
rect 18408 1776 18426 1840
rect 18490 1776 18508 1840
rect 18572 1776 18590 1840
rect 18654 1776 18660 1840
rect 17675 1754 18660 1776
rect 17675 1690 17681 1754
rect 17745 1690 17764 1754
rect 17828 1690 17847 1754
rect 17911 1690 17930 1754
rect 17994 1690 18013 1754
rect 18077 1690 18096 1754
rect 18160 1690 18179 1754
rect 18243 1690 18262 1754
rect 18326 1690 18344 1754
rect 18408 1690 18426 1754
rect 18490 1690 18508 1754
rect 18572 1690 18590 1754
rect 18654 1690 18660 1754
rect 17675 1668 18660 1690
rect 17675 1604 17681 1668
rect 17745 1604 17764 1668
rect 17828 1604 17847 1668
rect 17911 1604 17930 1668
rect 17994 1604 18013 1668
rect 18077 1604 18096 1668
rect 18160 1604 18179 1668
rect 18243 1604 18262 1668
rect 18326 1604 18344 1668
rect 18408 1604 18426 1668
rect 18490 1604 18508 1668
rect 18572 1604 18590 1668
rect 18654 1604 18660 1668
rect 17675 1582 18660 1604
rect 17675 1518 17681 1582
rect 17745 1518 17764 1582
rect 17828 1518 17847 1582
rect 17911 1518 17930 1582
rect 17994 1518 18013 1582
rect 18077 1518 18096 1582
rect 18160 1518 18179 1582
rect 18243 1518 18262 1582
rect 18326 1518 18344 1582
rect 18408 1518 18426 1582
rect 18490 1518 18508 1582
rect 18572 1518 18590 1582
rect 18654 1518 18660 1582
rect 17675 1514 18660 1518
tri 18839 1860 18885 1906 se
rect 18885 1860 19227 2109
rect 20734 2097 21132 2121
rect 20734 2041 20743 2097
rect 20799 2041 20825 2097
rect 20881 2041 20907 2097
rect 20963 2041 20989 2097
rect 21045 2041 21071 2097
rect 21127 2041 21132 2097
rect 20734 2036 21132 2041
rect 18839 1122 19227 1860
rect 18839 1076 18848 1122
rect 18904 1076 18929 1122
rect 18985 1076 19010 1122
rect 19066 1076 19227 1122
rect 17486 1045 17552 1050
rect 17486 989 17491 1045
rect 17547 989 17552 1045
rect 17486 965 17552 989
rect 17486 909 17491 965
rect 17547 909 17552 965
rect 17486 904 17552 909
rect 18839 1012 18842 1076
rect 18906 1012 18922 1076
rect 18986 1012 19002 1076
rect 19066 1012 19082 1076
rect 19146 1012 19162 1076
rect 19226 1012 19227 1076
rect 18839 996 19227 1012
rect 18839 991 18848 996
rect 18904 991 18929 996
rect 18985 991 19010 996
rect 19066 991 19227 996
rect 18839 927 18842 991
rect 18906 927 18922 991
rect 18986 927 19002 991
rect 19066 927 19082 991
rect 19146 927 19162 991
rect 19226 927 19227 991
rect 18839 906 19227 927
rect 18839 842 18842 906
rect 18906 842 18922 906
rect 18986 842 19002 906
rect 19066 842 19082 906
rect 19146 842 19162 906
rect 19226 842 19227 906
rect 18839 821 19227 842
rect 18839 757 18842 821
rect 18906 757 18922 821
rect 18986 757 19002 821
rect 19066 757 19082 821
rect 19146 757 19162 821
rect 19226 757 19227 821
rect 18839 736 19227 757
rect 18839 672 18842 736
rect 18906 672 18922 736
rect 18986 672 19002 736
rect 19066 672 19082 736
rect 19146 672 19162 736
rect 19226 672 19227 736
rect 18839 651 19227 672
rect 24857 718 24939 723
rect 24857 662 24875 718
rect 24931 662 24939 718
rect 18839 587 18842 651
rect 18906 587 18922 651
rect 18986 587 19002 651
rect 19066 587 19082 651
rect 19146 587 19162 651
rect 19226 587 19227 651
rect 18839 566 19227 587
rect 18839 502 18842 566
rect 18906 502 18922 566
rect 18986 502 19002 566
rect 19066 502 19082 566
rect 19146 502 19162 566
rect 19226 502 19227 566
rect 18839 481 19227 502
rect 18839 417 18842 481
rect 18906 417 18922 481
rect 18986 417 19002 481
rect 19066 417 19082 481
rect 19146 417 19162 481
rect 19226 417 19227 481
rect 18839 396 19227 417
rect 18839 332 18842 396
rect 18906 332 18922 396
rect 18986 332 19002 396
rect 19066 332 19082 396
rect 19146 332 19162 396
rect 19226 332 19227 396
rect 18839 311 19227 332
rect 18839 247 18842 311
rect 18906 247 18922 311
rect 18986 247 19002 311
rect 19066 247 19082 311
rect 19146 247 19162 311
rect 19226 247 19227 311
rect 18839 225 19227 247
rect 18839 161 18842 225
rect 18906 161 18922 225
rect 18986 161 19002 225
rect 19066 161 19082 225
rect 19146 161 19162 225
rect 19226 161 19227 225
rect 18839 154 19227 161
rect 24496 650 24562 655
rect 24496 594 24501 650
rect 24557 594 24562 650
rect 24496 570 24562 594
rect 24496 514 24501 570
rect 24557 514 24562 570
tri 17426 83 17441 98 sw
rect 17326 78 17472 83
rect 17326 22 17331 78
rect 17387 22 17411 78
rect 17467 22 17472 78
rect 17326 17 17472 22
rect 13243 -13 13825 -8
rect 13243 -69 13248 -13
rect 13304 -69 13352 -13
rect 13408 -69 13455 -13
rect 13511 -69 13558 -13
rect 13614 -69 13661 -13
rect 13717 -69 13764 -13
rect 13820 -69 13825 -13
rect 13243 -113 13825 -69
rect 13243 -169 13248 -113
rect 13304 -169 13352 -113
rect 13408 -169 13455 -113
rect 13511 -169 13558 -113
rect 13614 -169 13661 -113
rect 13717 -169 13764 -113
rect 13820 -169 13825 -113
rect 13243 -174 13825 -169
tri 7852 -409 7998 -263 nw
tri 7596 -452 7639 -409 se
rect 7639 -452 7809 -409
tri 7809 -452 7852 -409 nw
rect 634 -1103 766 -1096
rect 634 -1167 668 -1103
rect 732 -1167 766 -1103
rect 634 -1190 766 -1167
rect 634 -1254 668 -1190
rect 732 -1254 766 -1190
rect 634 -1277 766 -1254
rect 634 -1341 668 -1277
rect 732 -1341 766 -1277
rect 634 -1364 766 -1341
rect 634 -1428 668 -1364
rect 732 -1428 766 -1364
rect 634 -1451 766 -1428
rect 634 -1515 668 -1451
rect 732 -1515 766 -1451
rect 634 -1539 766 -1515
rect 634 -1603 668 -1539
rect 732 -1603 766 -1539
rect 634 -1627 766 -1603
rect 634 -1691 668 -1627
rect 732 -1691 766 -1627
rect 634 -1715 766 -1691
rect 634 -1779 668 -1715
rect 732 -1779 766 -1715
rect 634 -4288 766 -1779
rect 7596 -1105 7784 -452
tri 7784 -477 7809 -452 nw
rect 7596 -1169 7598 -1105
rect 7662 -1169 7718 -1105
rect 7782 -1169 7784 -1105
rect 7596 -1192 7784 -1169
rect 7596 -1256 7598 -1192
rect 7662 -1256 7718 -1192
rect 7782 -1256 7784 -1192
rect 7596 -1279 7784 -1256
rect 7596 -1343 7598 -1279
rect 7662 -1343 7718 -1279
rect 7782 -1343 7784 -1279
rect 7596 -1366 7784 -1343
rect 7596 -1430 7598 -1366
rect 7662 -1430 7718 -1366
rect 7782 -1430 7784 -1366
rect 7596 -1453 7784 -1430
rect 7596 -1517 7598 -1453
rect 7662 -1517 7718 -1453
rect 7782 -1517 7784 -1453
rect 7596 -1540 7784 -1517
rect 7596 -1604 7598 -1540
rect 7662 -1604 7718 -1540
rect 7782 -1604 7784 -1540
rect 7596 -1627 7784 -1604
rect 7596 -1691 7598 -1627
rect 7662 -1691 7718 -1627
rect 7782 -1691 7784 -1627
rect 7596 -1715 7784 -1691
rect 7596 -1779 7598 -1715
rect 7662 -1779 7718 -1715
rect 7782 -1779 7784 -1715
rect 7596 -1787 7784 -1779
rect 24496 -1713 24562 514
rect 24857 638 24939 662
rect 24857 582 24875 638
rect 24931 582 24939 638
rect 24857 -132 24939 582
rect 24857 -196 24866 -132
rect 24930 -196 24939 -132
rect 24857 -219 24939 -196
rect 24857 -283 24866 -219
rect 24930 -283 24939 -219
rect 24857 -306 24939 -283
rect 24857 -370 24866 -306
rect 24930 -370 24939 -306
rect 24857 -394 24939 -370
rect 24857 -458 24866 -394
rect 24930 -458 24939 -394
rect 24857 -482 24939 -458
rect 24857 -546 24866 -482
rect 24930 -546 24939 -482
rect 24857 -570 24939 -546
rect 24857 -634 24866 -570
rect 24930 -634 24939 -570
rect 24857 -658 24939 -634
rect 24857 -722 24866 -658
rect 24930 -722 24939 -658
rect 24857 -746 24939 -722
rect 24857 -810 24866 -746
rect 24930 -810 24939 -746
rect 24857 -816 24939 -810
rect 24496 -1769 24501 -1713
rect 24557 -1769 24562 -1713
rect 24496 -1793 24562 -1769
rect 24496 -1849 24501 -1793
rect 24557 -1849 24562 -1793
rect 24496 -1854 24562 -1849
rect 634 -4344 666 -4288
rect 722 -4344 766 -4288
rect 634 -4368 766 -4344
rect 634 -4424 666 -4368
rect 722 -4424 766 -4368
rect 634 -4429 766 -4424
rect 23354 -2005 23420 -2000
rect 23354 -2061 23359 -2005
rect 23415 -2061 23420 -2005
rect 23354 -2085 23420 -2061
rect 23354 -2141 23359 -2085
rect 23415 -2141 23420 -2085
rect 23354 -4492 23420 -2141
rect 633 -7756 765 -4518
rect 23354 -4556 23355 -4492
rect 23419 -4556 23420 -4492
rect 23354 -4579 23420 -4556
rect 23354 -4643 23355 -4579
rect 23419 -4643 23420 -4579
rect 23354 -4666 23420 -4643
rect 23354 -4730 23355 -4666
rect 23419 -4730 23420 -4666
rect 23354 -4753 23420 -4730
rect 23354 -4817 23355 -4753
rect 23419 -4817 23420 -4753
rect 23354 -4841 23420 -4817
rect 23354 -4905 23355 -4841
rect 23419 -4905 23420 -4841
rect 23354 -4929 23420 -4905
rect 23354 -4993 23355 -4929
rect 23419 -4993 23420 -4929
rect 23354 -5017 23420 -4993
rect 23354 -5081 23355 -5017
rect 23419 -5081 23420 -5017
rect 23354 -5105 23420 -5081
rect 23354 -5169 23355 -5105
rect 23419 -5169 23420 -5105
rect 23354 -5174 23420 -5169
rect 23355 -5175 23419 -5174
<< via3 >>
rect 20740 5440 20804 5504
rect 20820 5440 20884 5504
rect 20900 5440 20964 5504
rect 20980 5440 21044 5504
rect 21060 5440 21124 5504
rect 20740 5354 20804 5418
rect 20820 5354 20884 5418
rect 20900 5354 20964 5418
rect 20980 5354 21044 5418
rect 21060 5354 21124 5418
rect 20740 5268 20804 5332
rect 20820 5268 20884 5332
rect 20900 5268 20964 5332
rect 20980 5268 21044 5332
rect 21060 5268 21124 5332
rect 20740 5182 20804 5246
rect 20820 5182 20884 5246
rect 20900 5182 20964 5246
rect 20980 5182 21044 5246
rect 21060 5182 21124 5246
rect 20740 5096 20804 5160
rect 20820 5096 20884 5160
rect 20900 5096 20964 5160
rect 20980 5096 21044 5160
rect 21060 5096 21124 5160
rect 20740 5010 20804 5074
rect 20820 5010 20884 5074
rect 20900 5010 20964 5074
rect 20980 5010 21044 5074
rect 21060 5010 21124 5074
rect 20740 4924 20804 4988
rect 20820 4924 20884 4988
rect 20900 4924 20964 4988
rect 20980 4924 21044 4988
rect 21060 4924 21124 4988
rect 20740 4838 20804 4902
rect 20820 4838 20884 4902
rect 20900 4838 20964 4902
rect 20980 4838 21044 4902
rect 21060 4838 21124 4902
rect 20740 4751 20804 4815
rect 20820 4751 20884 4815
rect 20900 4751 20964 4815
rect 20980 4751 21044 4815
rect 21060 4751 21124 4815
rect 20740 4664 20804 4728
rect 20820 4664 20884 4728
rect 20900 4664 20964 4728
rect 20980 4664 21044 4728
rect 21060 4664 21124 4728
rect 6447 2985 6511 3049
rect 6540 2985 6604 3049
rect 6632 2985 6696 3049
rect 6724 2985 6788 3049
rect 6816 2985 6880 3049
rect 6908 2985 6972 3049
rect 7000 2985 7064 3049
rect 6447 2899 6511 2963
rect 6540 2899 6604 2963
rect 6632 2899 6696 2963
rect 6724 2899 6788 2963
rect 6816 2899 6880 2963
rect 6908 2899 6972 2963
rect 7000 2899 7064 2963
rect 6447 2813 6511 2877
rect 6540 2813 6604 2877
rect 6632 2813 6696 2877
rect 6724 2813 6788 2877
rect 6816 2813 6880 2877
rect 6908 2813 6972 2877
rect 7000 2813 7064 2877
rect 6447 2727 6511 2791
rect 6540 2727 6604 2791
rect 6632 2727 6696 2791
rect 6724 2727 6788 2791
rect 6816 2727 6880 2791
rect 6908 2727 6972 2791
rect 7000 2727 7064 2791
rect 6447 2641 6511 2705
rect 6540 2641 6604 2705
rect 6632 2641 6696 2705
rect 6724 2641 6788 2705
rect 6816 2641 6880 2705
rect 6908 2641 6972 2705
rect 7000 2641 7064 2705
rect 6447 2555 6511 2619
rect 6540 2555 6604 2619
rect 6632 2555 6696 2619
rect 6724 2555 6788 2619
rect 6816 2555 6880 2619
rect 6908 2555 6972 2619
rect 7000 2555 7064 2619
rect 6447 2469 6511 2533
rect 6540 2469 6604 2533
rect 6632 2469 6696 2533
rect 6724 2469 6788 2533
rect 6816 2469 6880 2533
rect 6908 2469 6972 2533
rect 7000 2469 7064 2533
rect 7875 2985 7939 3049
rect 7969 2985 8033 3049
rect 8062 2985 8126 3049
rect 8155 2985 8219 3049
rect 8248 2985 8312 3049
rect 8341 2985 8405 3049
rect 8434 2985 8498 3049
rect 7875 2899 7939 2963
rect 7969 2899 8033 2963
rect 8062 2899 8126 2963
rect 8155 2899 8219 2963
rect 8248 2899 8312 2963
rect 8341 2899 8405 2963
rect 8434 2899 8498 2963
rect 7875 2813 7939 2877
rect 7969 2813 8033 2877
rect 8062 2813 8126 2877
rect 8155 2813 8219 2877
rect 8248 2813 8312 2877
rect 8341 2813 8405 2877
rect 8434 2813 8498 2877
rect 7875 2727 7939 2791
rect 7969 2727 8033 2791
rect 8062 2727 8126 2791
rect 8155 2727 8219 2791
rect 8248 2727 8312 2791
rect 8341 2727 8405 2791
rect 8434 2727 8498 2791
rect 7875 2641 7939 2705
rect 7969 2641 8033 2705
rect 8062 2641 8126 2705
rect 8155 2641 8219 2705
rect 8248 2641 8312 2705
rect 8341 2641 8405 2705
rect 8434 2641 8498 2705
rect 7875 2555 7939 2619
rect 7969 2555 8033 2619
rect 8062 2555 8126 2619
rect 8155 2555 8219 2619
rect 8248 2555 8312 2619
rect 8341 2555 8405 2619
rect 8434 2555 8498 2619
rect 7875 2469 7939 2533
rect 7969 2469 8033 2533
rect 8062 2469 8126 2533
rect 8155 2469 8219 2533
rect 8248 2469 8312 2533
rect 8341 2469 8405 2533
rect 8434 2469 8498 2533
rect 15885 2034 15949 2098
rect 15978 2034 16042 2098
rect 16070 2034 16134 2098
rect 16162 2034 16226 2098
rect 16254 2034 16318 2098
rect 16346 2034 16410 2098
rect 16438 2034 16502 2098
rect 15885 1948 15949 2012
rect 15978 1948 16042 2012
rect 16070 1948 16134 2012
rect 16162 1948 16226 2012
rect 16254 1948 16318 2012
rect 16346 1948 16410 2012
rect 16438 1948 16502 2012
rect 15885 1862 15949 1926
rect 15978 1862 16042 1926
rect 16070 1862 16134 1926
rect 16162 1862 16226 1926
rect 16254 1862 16318 1926
rect 16346 1862 16410 1926
rect 16438 1862 16502 1926
rect 15885 1776 15949 1840
rect 15978 1776 16042 1840
rect 16070 1776 16134 1840
rect 16162 1776 16226 1840
rect 16254 1776 16318 1840
rect 16346 1776 16410 1840
rect 16438 1776 16502 1840
rect 15885 1690 15949 1754
rect 15978 1690 16042 1754
rect 16070 1690 16134 1754
rect 16162 1690 16226 1754
rect 16254 1690 16318 1754
rect 16346 1690 16410 1754
rect 16438 1690 16502 1754
rect 15885 1604 15949 1668
rect 15978 1604 16042 1668
rect 16070 1604 16134 1668
rect 16162 1604 16226 1668
rect 16254 1604 16318 1668
rect 16346 1604 16410 1668
rect 16438 1604 16502 1668
rect 15885 1518 15949 1582
rect 15978 1518 16042 1582
rect 16070 1518 16134 1582
rect 16162 1518 16226 1582
rect 16254 1518 16318 1582
rect 16346 1518 16410 1582
rect 16438 1518 16502 1582
rect 17681 2034 17745 2098
rect 17764 2034 17828 2098
rect 17847 2034 17911 2098
rect 17930 2034 17994 2098
rect 18013 2034 18077 2098
rect 18096 2034 18160 2098
rect 18179 2034 18243 2098
rect 18262 2034 18326 2098
rect 18344 2034 18408 2098
rect 18426 2034 18490 2098
rect 18508 2034 18572 2098
rect 18590 2034 18654 2098
rect 17681 1948 17745 2012
rect 17764 1948 17828 2012
rect 17847 1948 17911 2012
rect 17930 1948 17994 2012
rect 18013 1948 18077 2012
rect 18096 1948 18160 2012
rect 18179 1948 18243 2012
rect 18262 1948 18326 2012
rect 18344 1948 18408 2012
rect 18426 1948 18490 2012
rect 18508 1948 18572 2012
rect 18590 1948 18654 2012
rect 17681 1862 17745 1926
rect 17764 1862 17828 1926
rect 17847 1862 17911 1926
rect 17930 1862 17994 1926
rect 18013 1862 18077 1926
rect 18096 1862 18160 1926
rect 18179 1862 18243 1926
rect 18262 1862 18326 1926
rect 18344 1862 18408 1926
rect 18426 1862 18490 1926
rect 18508 1862 18572 1926
rect 18590 1862 18654 1926
rect 17681 1776 17745 1840
rect 17764 1776 17828 1840
rect 17847 1776 17911 1840
rect 17930 1776 17994 1840
rect 18013 1776 18077 1840
rect 18096 1776 18160 1840
rect 18179 1776 18243 1840
rect 18262 1776 18326 1840
rect 18344 1776 18408 1840
rect 18426 1776 18490 1840
rect 18508 1776 18572 1840
rect 18590 1776 18654 1840
rect 17681 1690 17745 1754
rect 17764 1690 17828 1754
rect 17847 1690 17911 1754
rect 17930 1690 17994 1754
rect 18013 1690 18077 1754
rect 18096 1690 18160 1754
rect 18179 1690 18243 1754
rect 18262 1690 18326 1754
rect 18344 1690 18408 1754
rect 18426 1690 18490 1754
rect 18508 1690 18572 1754
rect 18590 1690 18654 1754
rect 17681 1604 17745 1668
rect 17764 1604 17828 1668
rect 17847 1604 17911 1668
rect 17930 1604 17994 1668
rect 18013 1604 18077 1668
rect 18096 1604 18160 1668
rect 18179 1604 18243 1668
rect 18262 1604 18326 1668
rect 18344 1604 18408 1668
rect 18426 1604 18490 1668
rect 18508 1604 18572 1668
rect 18590 1604 18654 1668
rect 17681 1518 17745 1582
rect 17764 1518 17828 1582
rect 17847 1518 17911 1582
rect 17930 1518 17994 1582
rect 18013 1518 18077 1582
rect 18096 1518 18160 1582
rect 18179 1518 18243 1582
rect 18262 1518 18326 1582
rect 18344 1518 18408 1582
rect 18426 1518 18490 1582
rect 18508 1518 18572 1582
rect 18590 1518 18654 1582
rect 18842 1066 18848 1076
rect 18848 1066 18904 1076
rect 18904 1066 18906 1076
rect 18842 1012 18906 1066
rect 18922 1066 18929 1076
rect 18929 1066 18985 1076
rect 18985 1066 18986 1076
rect 18922 1012 18986 1066
rect 19002 1066 19010 1076
rect 19010 1066 19066 1076
rect 19002 1012 19066 1066
rect 19082 1012 19146 1076
rect 19162 1012 19226 1076
rect 18842 940 18848 991
rect 18848 940 18904 991
rect 18904 940 18906 991
rect 18842 927 18906 940
rect 18922 940 18929 991
rect 18929 940 18985 991
rect 18985 940 18986 991
rect 18922 927 18986 940
rect 19002 940 19010 991
rect 19010 940 19066 991
rect 19002 927 19066 940
rect 19082 927 19146 991
rect 19162 927 19226 991
rect 18842 842 18906 906
rect 18922 842 18986 906
rect 19002 842 19066 906
rect 19082 842 19146 906
rect 19162 842 19226 906
rect 18842 757 18906 821
rect 18922 757 18986 821
rect 19002 757 19066 821
rect 19082 757 19146 821
rect 19162 757 19226 821
rect 18842 672 18906 736
rect 18922 672 18986 736
rect 19002 672 19066 736
rect 19082 672 19146 736
rect 19162 672 19226 736
rect 18842 587 18906 651
rect 18922 587 18986 651
rect 19002 587 19066 651
rect 19082 587 19146 651
rect 19162 587 19226 651
rect 18842 502 18906 566
rect 18922 502 18986 566
rect 19002 502 19066 566
rect 19082 502 19146 566
rect 19162 502 19226 566
rect 18842 417 18906 481
rect 18922 417 18986 481
rect 19002 417 19066 481
rect 19082 417 19146 481
rect 19162 417 19226 481
rect 18842 332 18906 396
rect 18922 332 18986 396
rect 19002 332 19066 396
rect 19082 332 19146 396
rect 19162 332 19226 396
rect 18842 247 18906 311
rect 18922 247 18986 311
rect 19002 247 19066 311
rect 19082 247 19146 311
rect 19162 247 19226 311
rect 18842 161 18906 225
rect 18922 161 18986 225
rect 19002 161 19066 225
rect 19082 161 19146 225
rect 19162 161 19226 225
rect 668 -1167 732 -1103
rect 668 -1254 732 -1190
rect 668 -1341 732 -1277
rect 668 -1428 732 -1364
rect 668 -1515 732 -1451
rect 668 -1603 732 -1539
rect 668 -1691 732 -1627
rect 668 -1779 732 -1715
rect 7598 -1169 7662 -1105
rect 7718 -1169 7782 -1105
rect 7598 -1256 7662 -1192
rect 7718 -1256 7782 -1192
rect 7598 -1343 7662 -1279
rect 7718 -1343 7782 -1279
rect 7598 -1430 7662 -1366
rect 7718 -1430 7782 -1366
rect 7598 -1517 7662 -1453
rect 7718 -1517 7782 -1453
rect 7598 -1604 7662 -1540
rect 7718 -1604 7782 -1540
rect 7598 -1691 7662 -1627
rect 7718 -1691 7782 -1627
rect 7598 -1779 7662 -1715
rect 7718 -1779 7782 -1715
rect 24866 -196 24930 -132
rect 24866 -283 24930 -219
rect 24866 -370 24930 -306
rect 24866 -458 24930 -394
rect 24866 -546 24930 -482
rect 24866 -634 24930 -570
rect 24866 -722 24930 -658
rect 24866 -810 24930 -746
rect 23355 -4556 23419 -4492
rect 23355 -4643 23419 -4579
rect 23355 -4730 23419 -4666
rect 23355 -4817 23419 -4753
rect 23355 -4905 23419 -4841
rect 23355 -4993 23419 -4929
rect 23355 -5081 23419 -5017
rect 23355 -5169 23419 -5105
<< metal4 >>
rect 20738 5504 21126 5505
rect 20738 5440 20740 5504
rect 20804 5440 20820 5504
rect 20884 5440 20900 5504
rect 20964 5440 20980 5504
rect 21044 5440 21060 5504
rect 21124 5440 21126 5504
rect 20738 5418 21126 5440
rect 20738 5354 20740 5418
rect 20804 5354 20820 5418
rect 20884 5354 20900 5418
rect 20964 5354 20980 5418
rect 21044 5354 21060 5418
rect 21124 5354 21126 5418
rect 20738 5332 21126 5354
rect 20738 5268 20740 5332
rect 20804 5268 20820 5332
rect 20884 5268 20900 5332
rect 20964 5268 20980 5332
rect 21044 5268 21060 5332
rect 21124 5268 21126 5332
rect 20738 5246 21126 5268
rect 20738 5182 20740 5246
rect 20804 5182 20820 5246
rect 20884 5182 20900 5246
rect 20964 5182 20980 5246
rect 21044 5182 21060 5246
rect 21124 5182 21126 5246
rect 20738 5160 21126 5182
rect 20738 5096 20740 5160
rect 20804 5096 20820 5160
rect 20884 5096 20900 5160
rect 20964 5096 20980 5160
rect 21044 5096 21060 5160
rect 21124 5096 21126 5160
rect 20738 5074 21126 5096
rect 20738 5010 20740 5074
rect 20804 5010 20820 5074
rect 20884 5010 20900 5074
rect 20964 5010 20980 5074
rect 21044 5010 21060 5074
rect 21124 5010 21126 5074
rect 20738 4988 21126 5010
rect 20738 4924 20740 4988
rect 20804 4924 20820 4988
rect 20884 4924 20900 4988
rect 20964 4924 20980 4988
rect 21044 4924 21060 4988
rect 21124 4924 21126 4988
rect 20738 4902 21126 4924
rect 20738 4838 20740 4902
rect 20804 4838 20820 4902
rect 20884 4838 20900 4902
rect 20964 4838 20980 4902
rect 21044 4838 21060 4902
rect 21124 4838 21126 4902
rect 20738 4815 21126 4838
rect 20738 4751 20740 4815
rect 20804 4751 20820 4815
rect 20884 4751 20900 4815
rect 20964 4751 20980 4815
rect 21044 4751 21060 4815
rect 21124 4751 21126 4815
rect 20738 4728 21126 4751
rect 20738 4664 20740 4728
rect 20804 4664 20820 4728
rect 20884 4664 20900 4728
rect 20964 4664 20980 4728
rect 21044 4664 21060 4728
rect 21124 4664 21126 4728
rect 20738 4663 21126 4664
rect 6446 3049 8499 3054
rect 6446 2985 6447 3049
rect 6511 2985 6540 3049
rect 6604 2985 6632 3049
rect 6696 2985 6724 3049
rect 6788 2985 6816 3049
rect 6880 2985 6908 3049
rect 6972 2985 7000 3049
rect 7064 2985 7875 3049
rect 7939 2985 7969 3049
rect 8033 2985 8062 3049
rect 8126 2985 8155 3049
rect 8219 2985 8248 3049
rect 8312 2985 8341 3049
rect 8405 2985 8434 3049
rect 8498 2985 8499 3049
rect 6446 2963 8499 2985
rect 6446 2899 6447 2963
rect 6511 2899 6540 2963
rect 6604 2899 6632 2963
rect 6696 2899 6724 2963
rect 6788 2899 6816 2963
rect 6880 2899 6908 2963
rect 6972 2899 7000 2963
rect 7064 2899 7875 2963
rect 7939 2899 7969 2963
rect 8033 2899 8062 2963
rect 8126 2899 8155 2963
rect 8219 2899 8248 2963
rect 8312 2899 8341 2963
rect 8405 2899 8434 2963
rect 8498 2899 8499 2963
rect 6446 2877 8499 2899
rect 6446 2813 6447 2877
rect 6511 2813 6540 2877
rect 6604 2813 6632 2877
rect 6696 2813 6724 2877
rect 6788 2813 6816 2877
rect 6880 2813 6908 2877
rect 6972 2813 7000 2877
rect 7064 2813 7875 2877
rect 7939 2813 7969 2877
rect 8033 2813 8062 2877
rect 8126 2813 8155 2877
rect 8219 2813 8248 2877
rect 8312 2813 8341 2877
rect 8405 2813 8434 2877
rect 8498 2813 8499 2877
rect 6446 2791 8499 2813
rect 6446 2727 6447 2791
rect 6511 2727 6540 2791
rect 6604 2727 6632 2791
rect 6696 2727 6724 2791
rect 6788 2727 6816 2791
rect 6880 2727 6908 2791
rect 6972 2727 7000 2791
rect 7064 2727 7875 2791
rect 7939 2727 7969 2791
rect 8033 2727 8062 2791
rect 8126 2727 8155 2791
rect 8219 2727 8248 2791
rect 8312 2727 8341 2791
rect 8405 2727 8434 2791
rect 8498 2727 8499 2791
rect 6446 2705 8499 2727
rect 6446 2641 6447 2705
rect 6511 2641 6540 2705
rect 6604 2641 6632 2705
rect 6696 2641 6724 2705
rect 6788 2641 6816 2705
rect 6880 2641 6908 2705
rect 6972 2641 7000 2705
rect 7064 2641 7875 2705
rect 7939 2641 7969 2705
rect 8033 2641 8062 2705
rect 8126 2641 8155 2705
rect 8219 2641 8248 2705
rect 8312 2641 8341 2705
rect 8405 2641 8434 2705
rect 8498 2641 8499 2705
rect 6446 2619 8499 2641
rect 6446 2555 6447 2619
rect 6511 2555 6540 2619
rect 6604 2555 6632 2619
rect 6696 2555 6724 2619
rect 6788 2555 6816 2619
rect 6880 2555 6908 2619
rect 6972 2555 7000 2619
rect 7064 2555 7875 2619
rect 7939 2555 7969 2619
rect 8033 2555 8062 2619
rect 8126 2555 8155 2619
rect 8219 2555 8248 2619
rect 8312 2555 8341 2619
rect 8405 2555 8434 2619
rect 8498 2555 8499 2619
rect 6446 2533 8499 2555
rect 6446 2469 6447 2533
rect 6511 2469 6540 2533
rect 6604 2469 6632 2533
rect 6696 2469 6724 2533
rect 6788 2469 6816 2533
rect 6880 2469 6908 2533
rect 6972 2469 7000 2533
rect 7064 2469 7875 2533
rect 7939 2469 7969 2533
rect 8033 2469 8062 2533
rect 8126 2469 8155 2533
rect 8219 2469 8248 2533
rect 8312 2469 8341 2533
rect 8405 2469 8434 2533
rect 8498 2469 8499 2533
rect 6446 2464 8499 2469
rect 15884 2098 18655 2103
rect 15884 2034 15885 2098
rect 15949 2034 15978 2098
rect 16042 2034 16070 2098
rect 16134 2034 16162 2098
rect 16226 2034 16254 2098
rect 16318 2034 16346 2098
rect 16410 2034 16438 2098
rect 16502 2034 17681 2098
rect 17745 2034 17764 2098
rect 17828 2034 17847 2098
rect 17911 2034 17930 2098
rect 17994 2034 18013 2098
rect 18077 2034 18096 2098
rect 18160 2034 18179 2098
rect 18243 2034 18262 2098
rect 18326 2034 18344 2098
rect 18408 2034 18426 2098
rect 18490 2034 18508 2098
rect 18572 2034 18590 2098
rect 18654 2034 18655 2098
rect 15884 2012 18655 2034
rect 15884 1948 15885 2012
rect 15949 1948 15978 2012
rect 16042 1948 16070 2012
rect 16134 1948 16162 2012
rect 16226 1948 16254 2012
rect 16318 1948 16346 2012
rect 16410 1948 16438 2012
rect 16502 1948 17681 2012
rect 17745 1948 17764 2012
rect 17828 1948 17847 2012
rect 17911 1948 17930 2012
rect 17994 1948 18013 2012
rect 18077 1948 18096 2012
rect 18160 1948 18179 2012
rect 18243 1948 18262 2012
rect 18326 1948 18344 2012
rect 18408 1948 18426 2012
rect 18490 1948 18508 2012
rect 18572 1948 18590 2012
rect 18654 1948 18655 2012
rect 15884 1926 18655 1948
rect 15884 1862 15885 1926
rect 15949 1862 15978 1926
rect 16042 1862 16070 1926
rect 16134 1862 16162 1926
rect 16226 1862 16254 1926
rect 16318 1862 16346 1926
rect 16410 1862 16438 1926
rect 16502 1862 17681 1926
rect 17745 1862 17764 1926
rect 17828 1862 17847 1926
rect 17911 1862 17930 1926
rect 17994 1862 18013 1926
rect 18077 1862 18096 1926
rect 18160 1862 18179 1926
rect 18243 1862 18262 1926
rect 18326 1862 18344 1926
rect 18408 1862 18426 1926
rect 18490 1862 18508 1926
rect 18572 1862 18590 1926
rect 18654 1862 18655 1926
rect 15884 1840 18655 1862
rect 15884 1776 15885 1840
rect 15949 1776 15978 1840
rect 16042 1776 16070 1840
rect 16134 1776 16162 1840
rect 16226 1776 16254 1840
rect 16318 1776 16346 1840
rect 16410 1776 16438 1840
rect 16502 1776 17681 1840
rect 17745 1776 17764 1840
rect 17828 1776 17847 1840
rect 17911 1776 17930 1840
rect 17994 1776 18013 1840
rect 18077 1776 18096 1840
rect 18160 1776 18179 1840
rect 18243 1776 18262 1840
rect 18326 1776 18344 1840
rect 18408 1776 18426 1840
rect 18490 1776 18508 1840
rect 18572 1776 18590 1840
rect 18654 1776 18655 1840
rect 15884 1754 18655 1776
rect 15884 1690 15885 1754
rect 15949 1690 15978 1754
rect 16042 1690 16070 1754
rect 16134 1690 16162 1754
rect 16226 1690 16254 1754
rect 16318 1690 16346 1754
rect 16410 1690 16438 1754
rect 16502 1690 17681 1754
rect 17745 1690 17764 1754
rect 17828 1690 17847 1754
rect 17911 1690 17930 1754
rect 17994 1690 18013 1754
rect 18077 1690 18096 1754
rect 18160 1690 18179 1754
rect 18243 1690 18262 1754
rect 18326 1690 18344 1754
rect 18408 1690 18426 1754
rect 18490 1690 18508 1754
rect 18572 1690 18590 1754
rect 18654 1690 18655 1754
rect 15884 1668 18655 1690
rect 15884 1604 15885 1668
rect 15949 1604 15978 1668
rect 16042 1604 16070 1668
rect 16134 1604 16162 1668
rect 16226 1604 16254 1668
rect 16318 1604 16346 1668
rect 16410 1604 16438 1668
rect 16502 1604 17681 1668
rect 17745 1604 17764 1668
rect 17828 1604 17847 1668
rect 17911 1604 17930 1668
rect 17994 1604 18013 1668
rect 18077 1604 18096 1668
rect 18160 1604 18179 1668
rect 18243 1604 18262 1668
rect 18326 1604 18344 1668
rect 18408 1604 18426 1668
rect 18490 1604 18508 1668
rect 18572 1604 18590 1668
rect 18654 1604 18655 1668
rect 15884 1582 18655 1604
rect 15884 1518 15885 1582
rect 15949 1518 15978 1582
rect 16042 1518 16070 1582
rect 16134 1518 16162 1582
rect 16226 1518 16254 1582
rect 16318 1518 16346 1582
rect 16410 1518 16438 1582
rect 16502 1518 17681 1582
rect 17745 1518 17764 1582
rect 17828 1518 17847 1582
rect 17911 1518 17930 1582
rect 17994 1518 18013 1582
rect 18077 1518 18096 1582
rect 18160 1518 18179 1582
rect 18243 1518 18262 1582
rect 18326 1518 18344 1582
rect 18408 1518 18426 1582
rect 18490 1518 18508 1582
rect 18572 1518 18590 1582
rect 18654 1518 18655 1582
rect 15884 1513 18655 1518
rect 18841 1076 19227 1077
rect 18841 1012 18842 1076
rect 18906 1012 18922 1076
rect 18986 1012 19002 1076
rect 19066 1012 19082 1076
rect 19146 1012 19162 1076
rect 19226 1012 19227 1076
rect 18841 991 19227 1012
rect 18841 927 18842 991
rect 18906 927 18922 991
rect 18986 927 19002 991
rect 19066 927 19082 991
rect 19146 927 19162 991
rect 19226 927 19227 991
rect 18841 906 19227 927
rect 18841 842 18842 906
rect 18906 842 18922 906
rect 18986 842 19002 906
rect 19066 842 19082 906
rect 19146 842 19162 906
rect 19226 842 19227 906
rect 18841 821 19227 842
rect 18841 757 18842 821
rect 18906 757 18922 821
rect 18986 757 19002 821
rect 19066 757 19082 821
rect 19146 757 19162 821
rect 19226 757 19227 821
rect 18841 736 19227 757
rect 18841 672 18842 736
rect 18906 672 18922 736
rect 18986 672 19002 736
rect 19066 672 19082 736
rect 19146 672 19162 736
rect 19226 672 19227 736
rect 18841 651 19227 672
rect 18841 587 18842 651
rect 18906 587 18922 651
rect 18986 587 19002 651
rect 19066 587 19082 651
rect 19146 587 19162 651
rect 19226 587 19227 651
rect 18841 566 19227 587
rect 18841 502 18842 566
rect 18906 502 18922 566
rect 18986 502 19002 566
rect 19066 502 19082 566
rect 19146 502 19162 566
rect 19226 502 19227 566
rect 18841 481 19227 502
rect 18841 417 18842 481
rect 18906 417 18922 481
rect 18986 417 19002 481
rect 19066 417 19082 481
rect 19146 417 19162 481
rect 19226 417 19227 481
rect 18841 396 19227 417
rect 18841 332 18842 396
rect 18906 332 18922 396
rect 18986 332 19002 396
rect 19066 332 19082 396
rect 19146 332 19162 396
rect 19226 332 19227 396
rect 18841 311 19227 332
rect 18841 247 18842 311
rect 18906 247 18922 311
rect 18986 247 19002 311
rect 19066 247 19082 311
rect 19146 247 19162 311
rect 19226 247 19227 311
rect 18841 225 19227 247
rect 18841 161 18842 225
rect 18906 161 18922 225
rect 18986 161 19002 225
rect 19066 161 19082 225
rect 19146 161 19162 225
rect 19226 161 19227 225
rect 18841 160 19227 161
rect 24865 -132 24931 -131
rect 24865 -196 24866 -132
rect 24930 -196 24931 -132
rect 24865 -219 24931 -196
rect 24865 -283 24866 -219
rect 24930 -283 24931 -219
rect 24865 -306 24931 -283
rect 24865 -370 24866 -306
rect 24930 -370 24931 -306
rect 24865 -394 24931 -370
rect 24865 -458 24866 -394
rect 24930 -458 24931 -394
rect 24865 -482 24931 -458
rect 24865 -546 24866 -482
rect 24930 -546 24931 -482
rect 24865 -570 24931 -546
rect 24865 -634 24866 -570
rect 24930 -634 24931 -570
rect 24865 -658 24931 -634
rect 24865 -722 24866 -658
rect 24930 -722 24931 -658
rect 24865 -746 24931 -722
rect 24865 -810 24866 -746
rect 24930 -810 24931 -746
rect 24865 -811 24931 -810
rect 635 -1103 765 -1102
rect 635 -1167 668 -1103
rect 732 -1167 765 -1103
rect 635 -1190 765 -1167
rect 635 -1254 668 -1190
rect 732 -1254 765 -1190
rect 635 -1277 765 -1254
rect 635 -1341 668 -1277
rect 732 -1341 765 -1277
rect 635 -1364 765 -1341
rect 635 -1428 668 -1364
rect 732 -1428 765 -1364
rect 635 -1451 765 -1428
rect 635 -1515 668 -1451
rect 732 -1515 765 -1451
rect 635 -1539 765 -1515
rect 635 -1603 668 -1539
rect 732 -1603 765 -1539
rect 635 -1627 765 -1603
rect 635 -1691 668 -1627
rect 732 -1691 765 -1627
rect 635 -1715 765 -1691
rect 635 -1779 668 -1715
rect 732 -1779 765 -1715
rect 635 -1780 765 -1779
rect 7597 -1105 7783 -1104
rect 7597 -1169 7598 -1105
rect 7662 -1169 7718 -1105
rect 7782 -1169 7783 -1105
rect 7597 -1192 7783 -1169
rect 7597 -1256 7598 -1192
rect 7662 -1256 7718 -1192
rect 7782 -1256 7783 -1192
rect 7597 -1279 7783 -1256
rect 7597 -1343 7598 -1279
rect 7662 -1343 7718 -1279
rect 7782 -1343 7783 -1279
rect 7597 -1366 7783 -1343
rect 7597 -1430 7598 -1366
rect 7662 -1430 7718 -1366
rect 7782 -1430 7783 -1366
rect 7597 -1453 7783 -1430
rect 7597 -1517 7598 -1453
rect 7662 -1517 7718 -1453
rect 7782 -1517 7783 -1453
rect 7597 -1540 7783 -1517
rect 7597 -1604 7598 -1540
rect 7662 -1604 7718 -1540
rect 7782 -1604 7783 -1540
rect 7597 -1627 7783 -1604
rect 7597 -1691 7598 -1627
rect 7662 -1691 7718 -1627
rect 7782 -1691 7783 -1627
rect 7597 -1715 7783 -1691
rect 7597 -1779 7598 -1715
rect 7662 -1779 7718 -1715
rect 7782 -1779 7783 -1715
rect 7597 -1780 7783 -1779
rect 23354 -4492 23420 -4491
rect 23354 -4556 23355 -4492
rect 23419 -4556 23420 -4492
rect 23354 -4579 23420 -4556
rect 23354 -4643 23355 -4579
rect 23419 -4643 23420 -4579
rect 23354 -4666 23420 -4643
rect 23354 -4730 23355 -4666
rect 23419 -4730 23420 -4666
rect 23354 -4753 23420 -4730
rect 23354 -4817 23355 -4753
rect 23419 -4817 23420 -4753
rect 23354 -4841 23420 -4817
rect 23354 -4905 23355 -4841
rect 23419 -4905 23420 -4841
rect 23354 -4929 23420 -4905
rect 23354 -4993 23355 -4929
rect 23419 -4993 23420 -4929
rect 23354 -5017 23420 -4993
rect 23354 -5081 23355 -5017
rect 23419 -5081 23420 -5017
rect 23354 -5105 23420 -5081
rect 23354 -5169 23355 -5105
rect 23419 -5169 23420 -5105
rect 23354 -5170 23420 -5169
use sky130_fd_io__gpio_ovtv2_amux_ctl_logic_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_ctl_logic_i2c_fix_0
timestamp 1663361622
transform 1 0 0 0 1 0
box -1368 -8163 25113 3933
use sky130_fd_io__gpio_ovtv2_amux_switch  sky130_fd_io__gpio_ovtv2_amux_switch_0
timestamp 1663361622
transform 1 0 7103 0 1 7197
box -33 416 8691 910
use sky130_fd_io__gpio_ovtv2_amux_switch_1  sky130_fd_io__gpio_ovtv2_amux_switch_1_0
timestamp 1663361622
transform 1 0 627 0 1 3653
box -847 -2831 12071 1859
use sky130_fd_io__gpio_ovtv2_amux_switch_2  sky130_fd_io__gpio_ovtv2_amux_switch_2_0
timestamp 1663361622
transform -1 0 24533 0 1 3653
box -509 -2139 12071 2812
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1663361622
transform 0 -1 253 1 0 1314
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1663361622
transform 0 -1 -740 1 0 1314
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_2
timestamp 1663361622
transform 0 -1 253 1 0 2196
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_3
timestamp 1663361622
transform 0 -1 749 1 0 1314
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_4
timestamp 1663361622
transform 0 -1 749 1 0 2196
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_5
timestamp 1663361622
transform 0 -1 -740 1 0 2196
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_6
timestamp 1663361622
transform 0 -1 -243 1 0 1314
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_7
timestamp 1663361622
transform 0 -1 -243 1 0 2196
box 0 0 882 404
use sky130_fd_pr__nfet_01v8__example_5595914180834  sky130_fd_pr__nfet_01v8__example_5595914180834_0
timestamp 1663361622
transform 1 0 1333 0 1 21721
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_5595914180834  sky130_fd_pr__nfet_01v8__example_5595914180834_1
timestamp 1663361622
transform 1 0 1333 0 -1 21589
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808472  sky130_fd_pr__nfet_01v8__example_55959141808472_0
timestamp 1663361622
transform -1 0 24506 0 -1 3029
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808524  sky130_fd_pr__nfet_01v8__example_55959141808524_0
timestamp 1663361622
transform 1 0 24874 0 1 861
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808524  sky130_fd_pr__nfet_01v8__example_55959141808524_1
timestamp 1663361622
transform -1 0 24682 0 -1 945
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_0
timestamp 1663361622
transform 1 0 1289 0 -1 9699
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_1
timestamp 1663361622
transform 1 0 1732 0 -1 10495
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808469  sky130_fd_pr__pfet_01v8__example_55959141808469_0
timestamp 1663361622
transform 1 0 24386 0 1 2517
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808525  sky130_fd_pr__pfet_01v8__example_55959141808525_0
timestamp 1663361622
transform -1 0 6752 0 -1 2717
box -1 0 201 1
<< labels >>
flabel metal1 s 153 4288 442 4415 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal1 s 24702 4136 24991 4263 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal1 s 7531 3728 7598 3930 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew
flabel metal1 s 10368 1941 10394 1960 3 FreeSans 400 0 0 0 ANALOG_EN
port 3 nsew
flabel metal1 s 12736 2775 12754 2800 3 FreeSans 400 90 0 0 ANALOG_POL
port 4 nsew
flabel metal1 s 9221 2767 9239 2790 3 FreeSans 400 90 0 0 ANALOG_SEL
port 5 nsew
flabel metal1 s -294 -6430 -277 -6408 3 FreeSans 400 90 0 0 ENABLE_VDDA_H
port 6 nsew
flabel metal1 s -803 -5553 -780 -5527 3 FreeSans 400 90 0 0 ENABLE_VSWITCH_H
port 7 nsew
flabel metal1 s 12386 1917 12415 1943 3 FreeSans 400 0 0 0 OUT
port 8 nsew
flabel metal1 s 11939 1264 11976 1289 3 FreeSans 400 0 0 0 VCCD
port 9 nsew
flabel metal1 s 2255 3501 2320 3552 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal1 s 22292 2307 22323 2347 3 FreeSans 400 90 0 0 VDDIO_Q
port 10 nsew
flabel metal1 s 1144 22601 1183 22632 3 FreeSans 400 0 0 0 VSSIO
port 11 nsew
flabel metal1 s 7822 1038 7857 1068 3 FreeSans 400 0 0 0 VSWITCH
port 12 nsew
flabel metal1 s 23350 2706 23384 2741 3 FreeSans 400 90 0 0 PU_CSD_H
port 13 nsew
flabel metal1 s 707 -6388 744 -6358 3 FreeSans 400 0 0 0 VDDA
port 14 nsew
flabel metal1 s 6244 2465 6281 2495 3 FreeSans 400 0 0 0 VDDA
port 14 nsew
flabel metal1 s 15781 2472 15818 2502 3 FreeSans 400 0 0 0 VDDA
port 14 nsew
flabel metal1 s -1112 -6297 -1047 -6246 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal1 s 24734 755 24779 820 3 FreeSans 520 90 0 0 VSSA
port 1 nsew
flabel metal1 s -286 -4433 -251 -4403 3 FreeSans 400 0 0 0 VSWITCH
port 12 nsew
flabel metal1 s -613 -3123 -582 -3083 3 FreeSans 400 90 0 0 VDDIO_Q
port 10 nsew
flabel metal1 s 20866 2307 20897 2347 3 FreeSans 400 90 0 0 VDDIO_Q
port 10 nsew
flabel locali s 11396 8113 11463 8175 3 FreeSans 520 180 0 0 VPB_DRVR
port 15 nsew
flabel metal3 s 6602 2465 6856 3061 3 FreeSans 520 0 0 0 AMUXBUS_A
port 16 nsew
flabel metal3 s 16060 2200 16314 2796 3 FreeSans 520 0 0 0 AMUXBUS_B
port 17 nsew
flabel metal2 s 2419 10159 2471 10226 3 FreeSans 520 90 0 0 PGHS_H
port 18 nsew
flabel metal2 s 1854 22361 1921 22413 3 FreeSans 520 180 0 0 NGHS_H
port 19 nsew
flabel metal2 s -277 1014 -111 1114 3 FreeSans 520 180 0 0 PAD
port 20 nsew
flabel metal2 s 2258 5976 2305 6075 3 FreeSans 520 270 0 0 PUG_H[0]
port 21 nsew
flabel metal2 s 2340 5976 2387 6075 3 FreeSans 520 270 0 0 PUG_H[1]
port 22 nsew
flabel metal2 s 1307 1872 1347 1924 3 FreeSans 520 90 0 0 PD_CSD_H
port 23 nsew
flabel metal2 s 12187 4053 12233 4105 3 FreeSans 520 90 0 0 NGA_PAD_VPMP_H
port 24 nsew
flabel metal2 s 12930 4086 12968 4138 3 FreeSans 520 90 0 0 NGB_PAD_VPMP_H
port 25 nsew
flabel metal2 s 21019 1383 21042 1402 3 FreeSans 400 0 0 0 HLD_I_H_N
port 26 nsew
flabel metal2 s 22727 1293 22769 1325 3 FreeSans 400 0 0 0 VSSD
port 27 nsew
flabel metal2 s 11939 -1733 11976 -1708 3 FreeSans 400 0 0 0 VCCD
port 9 nsew
flabel comment s 2276 6036 2276 6036 0 FreeSans 400 90 0 0 PUG<0>
flabel comment s 2364 6036 2364 6036 0 FreeSans 400 90 0 0 PUG<1>
flabel comment s 7338 616 7338 616 0 FreeSans 2000 0 0 0 VSWITCH
flabel comment s 24733 972 24733 972 0 FreeSans 280 180 0 0 CONDIODE
<< properties >>
string GDS_END 31363332
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 30223726
<< end >>
