/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/ngspice/capacitors/sky130_fd_pr__model__cap_var.model.spice