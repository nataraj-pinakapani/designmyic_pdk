magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 268 163 459 203
rect 3 27 459 163
rect 28 -17 62 27
rect 268 21 459 27
<< locali >>
rect 17 425 255 483
rect 120 265 159 323
rect 387 299 442 493
rect 17 199 86 265
rect 120 199 285 265
rect 408 152 442 299
rect 387 83 442 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 21 357 255 391
rect 289 367 345 527
rect 21 299 86 357
rect 221 333 255 357
rect 221 299 353 333
rect 319 265 353 299
rect 319 199 374 265
rect 319 165 353 199
rect 20 131 353 165
rect 20 61 71 131
rect 105 17 171 97
rect 205 61 239 131
rect 273 17 349 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 120 199 285 265 6 A
port 1 nsew signal input
rlabel locali s 120 265 159 323 6 A
port 1 nsew signal input
rlabel locali s 17 425 255 483 6 B
port 2 nsew signal input
rlabel locali s 17 199 86 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 268 21 459 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 28 -17 62 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 3 27 459 163 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 268 163 459 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 387 83 442 152 6 X
port 8 nsew signal output
rlabel locali s 408 152 442 299 6 X
port 8 nsew signal output
rlabel locali s 387 299 442 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1016844
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1011774
<< end >>
