magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 98 157 1011 203
rect 1 21 1011 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 174 47 204 177
rect 258 47 288 177
rect 342 47 372 177
rect 426 47 456 177
rect 587 47 617 177
rect 671 47 701 177
rect 785 47 815 177
rect 903 47 933 177
<< scpmoshvt >>
rect 79 413 109 497
rect 174 297 204 497
rect 258 297 288 497
rect 342 297 372 497
rect 426 297 456 497
rect 587 297 617 497
rect 671 297 701 497
rect 785 297 815 497
rect 903 297 933 497
<< ndiff >>
rect 124 131 174 177
rect 27 101 79 131
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 174 131
rect 109 59 130 93
rect 164 59 174 93
rect 109 47 174 59
rect 204 101 258 177
rect 204 67 214 101
rect 248 67 258 101
rect 204 47 258 67
rect 288 94 342 177
rect 288 60 298 94
rect 332 60 342 94
rect 288 47 342 60
rect 372 101 426 177
rect 372 67 382 101
rect 416 67 426 101
rect 372 47 426 67
rect 456 89 587 177
rect 456 55 473 89
rect 507 55 587 89
rect 456 47 587 55
rect 617 47 671 177
rect 701 47 785 177
rect 815 47 903 177
rect 933 162 985 177
rect 933 128 943 162
rect 977 128 985 162
rect 933 94 985 128
rect 933 60 943 94
rect 977 60 985 94
rect 933 47 985 60
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 413 79 443
rect 109 485 174 497
rect 109 451 119 485
rect 153 451 174 485
rect 109 413 174 451
rect 124 297 174 413
rect 204 343 258 497
rect 204 309 214 343
rect 248 309 258 343
rect 204 297 258 309
rect 288 485 342 497
rect 288 451 298 485
rect 332 451 342 485
rect 288 297 342 451
rect 372 343 426 497
rect 372 309 382 343
rect 416 309 426 343
rect 372 297 426 309
rect 456 485 587 497
rect 456 451 466 485
rect 500 451 587 485
rect 456 297 587 451
rect 617 343 671 497
rect 617 309 627 343
rect 661 309 671 343
rect 617 297 671 309
rect 701 485 785 497
rect 701 451 711 485
rect 745 451 785 485
rect 701 297 785 451
rect 815 343 903 497
rect 815 309 859 343
rect 893 309 903 343
rect 815 297 903 309
rect 933 485 985 497
rect 933 451 943 485
rect 977 451 985 485
rect 933 297 985 451
<< ndiffc >>
rect 35 67 69 101
rect 130 59 164 93
rect 214 67 248 101
rect 298 60 332 94
rect 382 67 416 101
rect 473 55 507 89
rect 943 128 977 162
rect 943 60 977 94
<< pdiffc >>
rect 35 443 69 477
rect 119 451 153 485
rect 214 309 248 343
rect 298 451 332 485
rect 382 309 416 343
rect 466 451 500 485
rect 627 309 661 343
rect 711 451 745 485
rect 859 309 893 343
rect 943 451 977 485
<< poly >>
rect 79 497 109 523
rect 174 497 204 523
rect 258 497 288 523
rect 342 497 372 523
rect 426 497 456 523
rect 587 497 617 523
rect 671 497 701 523
rect 785 497 815 523
rect 903 497 933 523
rect 79 265 109 413
rect 174 265 204 297
rect 258 265 288 297
rect 342 265 372 297
rect 426 265 456 297
rect 587 265 617 297
rect 671 265 701 297
rect 785 265 815 297
rect 903 265 933 297
rect 78 249 132 265
rect 78 215 88 249
rect 122 215 132 249
rect 78 199 132 215
rect 174 249 490 265
rect 174 215 304 249
rect 338 215 372 249
rect 406 215 440 249
rect 474 215 490 249
rect 174 199 490 215
rect 563 249 617 265
rect 563 215 573 249
rect 607 215 617 249
rect 563 199 617 215
rect 659 249 713 265
rect 659 215 669 249
rect 703 215 713 249
rect 659 199 713 215
rect 785 249 839 265
rect 785 215 795 249
rect 829 215 839 249
rect 785 199 839 215
rect 903 249 990 265
rect 903 215 946 249
rect 980 215 990 249
rect 903 199 990 215
rect 79 131 109 199
rect 174 177 204 199
rect 258 177 288 199
rect 342 177 372 199
rect 426 177 456 199
rect 587 177 617 199
rect 671 177 701 199
rect 785 177 815 199
rect 903 177 933 199
rect 79 21 109 47
rect 174 21 204 47
rect 258 21 288 47
rect 342 21 372 47
rect 426 21 456 47
rect 587 21 617 47
rect 671 21 701 47
rect 785 21 815 47
rect 903 21 933 47
<< polycont >>
rect 88 215 122 249
rect 304 215 338 249
rect 372 215 406 249
rect 440 215 474 249
rect 573 215 607 249
rect 669 215 703 249
rect 795 215 829 249
rect 946 215 980 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 282 485 348 527
rect 282 451 298 485
rect 332 451 348 485
rect 450 485 516 527
rect 450 451 466 485
rect 500 451 516 485
rect 695 485 761 527
rect 695 451 711 485
rect 745 451 761 485
rect 927 485 993 527
rect 927 451 943 485
rect 977 451 993 485
rect 17 417 69 443
rect 17 383 980 417
rect 17 117 52 383
rect 88 249 158 327
rect 122 215 158 249
rect 88 153 158 215
rect 196 309 214 343
rect 248 309 382 343
rect 416 309 432 343
rect 476 309 627 343
rect 661 309 859 343
rect 893 309 909 343
rect 196 164 252 309
rect 476 249 510 309
rect 288 215 304 249
rect 338 215 372 249
rect 406 215 440 249
rect 474 215 510 249
rect 196 130 416 164
rect 17 101 69 117
rect 17 67 35 101
rect 214 101 248 130
rect 17 51 69 67
rect 114 93 180 94
rect 114 59 130 93
rect 164 59 180 93
rect 114 17 180 59
rect 382 101 416 130
rect 476 157 510 215
rect 573 249 617 265
rect 607 215 617 249
rect 573 199 617 215
rect 669 249 711 265
rect 703 215 711 249
rect 476 123 593 157
rect 669 151 711 215
rect 763 249 829 265
rect 763 215 795 249
rect 763 147 829 215
rect 946 249 980 383
rect 946 199 980 215
rect 214 51 248 67
rect 282 60 298 94
rect 332 60 348 94
rect 282 17 348 60
rect 559 94 593 123
rect 878 128 943 162
rect 977 128 993 162
rect 878 94 993 128
rect 382 51 416 67
rect 457 55 473 89
rect 507 55 523 89
rect 559 60 943 94
rect 977 60 993 94
rect 457 17 523 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 674 153 708 187 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 766 153 800 187 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 and4b_4
rlabel metal1 s 0 -48 1012 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 3081060
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3073382
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 25.300 0.000 
<< end >>
