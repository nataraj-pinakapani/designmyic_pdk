magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 22 22 22 23 6 C0
port 1 nsew
rlabel  s 22 21 22 22 6 C0
port 1 nsew
rlabel  s 22 19 22 20 6 C0
port 1 nsew
rlabel  s 22 18 22 19 6 C0
port 1 nsew
rlabel  s 22 17 22 18 6 C0
port 1 nsew
rlabel  s 22 15 22 16 6 C0
port 1 nsew
rlabel  s 22 14 22 15 6 C0
port 1 nsew
rlabel  s 22 13 22 14 6 C0
port 1 nsew
rlabel  s 22 12 22 13 6 C0
port 1 nsew
rlabel  s 22 10 22 11 6 C0
port 1 nsew
rlabel  s 22 9 22 10 6 C0
port 1 nsew
rlabel  s 22 8 22 9 6 C0
port 1 nsew
rlabel  s 22 7 22 8 6 C0
port 1 nsew
rlabel  s 22 5 22 6 6 C0
port 1 nsew
rlabel  s 22 4 22 5 6 C0
port 1 nsew
rlabel  s 22 3 22 4 6 C0
port 1 nsew
rlabel  s 22 2 22 2 6 C0
port 1 nsew
rlabel  s 22 0 22 1 8 C0
port 1 nsew
rlabel  s 17 22 22 22 6 C0
port 1 nsew
rlabel  s 17 20 22 21 6 C0
port 1 nsew
rlabel  s 17 19 22 19 6 C0
port 1 nsew
rlabel  s 17 18 22 18 6 C0
port 1 nsew
rlabel  s 17 16 22 17 6 C0
port 1 nsew
rlabel  s 17 15 22 15 6 C0
port 1 nsew
rlabel  s 17 14 22 14 6 C0
port 1 nsew
rlabel  s 17 13 22 13 6 C0
port 1 nsew
rlabel  s 17 10 22 10 6 C0
port 1 nsew
rlabel  s 17 9 22 9 6 C0
port 1 nsew
rlabel  s 17 8 22 8 6 C0
port 1 nsew
rlabel  s 17 6 22 7 6 C0
port 1 nsew
rlabel  s 17 5 22 5 6 C0
port 1 nsew
rlabel  s 17 4 22 4 6 C0
port 1 nsew
rlabel  s 17 2 22 3 6 C0
port 1 nsew
rlabel  s 17 1 22 2 6 C0
port 1 nsew
rlabel  s 11 22 11 23 6 C0
port 1 nsew
rlabel  s 11 21 11 22 6 C0
port 1 nsew
rlabel  s 11 19 11 20 6 C0
port 1 nsew
rlabel  s 11 18 11 19 6 C0
port 1 nsew
rlabel  s 11 17 11 18 6 C0
port 1 nsew
rlabel  s 11 15 11 16 6 C0
port 1 nsew
rlabel  s 11 14 11 15 6 C0
port 1 nsew
rlabel  s 11 13 11 14 6 C0
port 1 nsew
rlabel  s 11 12 11 13 6 C0
port 1 nsew
rlabel  s 11 10 11 11 6 C0
port 1 nsew
rlabel  s 11 9 11 10 6 C0
port 1 nsew
rlabel  s 11 8 11 9 6 C0
port 1 nsew
rlabel  s 11 7 11 8 6 C0
port 1 nsew
rlabel  s 11 5 11 6 6 C0
port 1 nsew
rlabel  s 11 4 11 5 6 C0
port 1 nsew
rlabel  s 11 3 11 4 6 C0
port 1 nsew
rlabel  s 11 2 11 2 6 C0
port 1 nsew
rlabel  s 11 0 11 1 8 C0
port 1 nsew
rlabel  s 6 22 16 22 6 C0
port 1 nsew
rlabel  s 6 20 16 21 6 C0
port 1 nsew
rlabel  s 6 19 16 19 6 C0
port 1 nsew
rlabel  s 6 18 16 18 6 C0
port 1 nsew
rlabel  s 6 16 16 17 6 C0
port 1 nsew
rlabel  s 6 15 16 15 6 C0
port 1 nsew
rlabel  s 6 14 16 14 6 C0
port 1 nsew
rlabel  s 6 13 16 13 6 C0
port 1 nsew
rlabel  s 6 10 16 10 6 C0
port 1 nsew
rlabel  s 6 9 16 9 6 C0
port 1 nsew
rlabel  s 6 8 16 8 6 C0
port 1 nsew
rlabel  s 6 6 16 7 6 C0
port 1 nsew
rlabel  s 6 5 16 5 6 C0
port 1 nsew
rlabel  s 6 4 16 4 6 C0
port 1 nsew
rlabel  s 6 2 16 3 6 C0
port 1 nsew
rlabel  s 6 1 16 2 6 C0
port 1 nsew
rlabel  s 0 23 22 23 6 C0
port 1 nsew
rlabel  s 0 22 0 23 4 C0
port 1 nsew
rlabel  s 0 22 5 22 6 C0
port 1 nsew
rlabel  s 0 21 0 22 4 C0
port 1 nsew
rlabel  s 0 20 5 21 6 C0
port 1 nsew
rlabel  s 0 19 0 20 4 C0
port 1 nsew
rlabel  s 0 19 5 19 6 C0
port 1 nsew
rlabel  s 0 18 0 19 4 C0
port 1 nsew
rlabel  s 0 18 5 18 6 C0
port 1 nsew
rlabel  s 0 17 0 18 4 C0
port 1 nsew
rlabel  s 0 16 5 17 6 C0
port 1 nsew
rlabel  s 0 15 0 16 4 C0
port 1 nsew
rlabel  s 0 15 5 15 6 C0
port 1 nsew
rlabel  s 0 14 0 15 4 C0
port 1 nsew
rlabel  s 0 14 5 14 6 C0
port 1 nsew
rlabel  s 0 13 0 14 4 C0
port 1 nsew
rlabel  s 0 13 5 13 6 C0
port 1 nsew
rlabel  s 0 12 0 13 4 C0
port 1 nsew
rlabel  s 0 11 22 12 6 C0
port 1 nsew
rlabel  s 0 10 0 11 4 C0
port 1 nsew
rlabel  s 0 10 5 10 6 C0
port 1 nsew
rlabel  s 0 9 0 10 4 C0
port 1 nsew
rlabel  s 0 9 5 9 6 C0
port 1 nsew
rlabel  s 0 8 0 9 4 C0
port 1 nsew
rlabel  s 0 8 5 8 6 C0
port 1 nsew
rlabel  s 0 7 0 8 4 C0
port 1 nsew
rlabel  s 0 6 5 7 6 C0
port 1 nsew
rlabel  s 0 5 0 6 4 C0
port 1 nsew
rlabel  s 0 5 5 5 6 C0
port 1 nsew
rlabel  s 0 4 0 5 4 C0
port 1 nsew
rlabel  s 0 4 5 4 6 C0
port 1 nsew
rlabel  s 0 3 0 4 4 C0
port 1 nsew
rlabel  s 0 2 5 3 6 C0
port 1 nsew
rlabel  s 0 2 0 2 4 C0
port 1 nsew
rlabel  s 0 1 5 2 6 C0
port 1 nsew
rlabel  s 0 0 0 1 2 C0
port 1 nsew
rlabel  s 0 0 22 0 8 C0
port 1 nsew
rlabel  s 17 21 17 22 6 C1
port 2 nsew
rlabel  s 17 20 17 21 6 C1
port 2 nsew
rlabel  s 17 19 17 20 6 C1
port 2 nsew
rlabel  s 17 17 17 18 6 C1
port 2 nsew
rlabel  s 17 16 17 17 6 C1
port 2 nsew
rlabel  s 17 15 17 16 6 C1
port 2 nsew
rlabel  s 17 13 17 14 6 C1
port 2 nsew
rlabel  s 17 12 17 13 6 C1
port 2 nsew
rlabel  s 17 10 17 11 6 C1
port 2 nsew
rlabel  s 17 9 17 10 6 C1
port 2 nsew
rlabel  s 17 7 17 8 6 C1
port 2 nsew
rlabel  s 17 6 17 7 6 C1
port 2 nsew
rlabel  s 17 5 17 6 6 C1
port 2 nsew
rlabel  s 17 3 17 4 6 C1
port 2 nsew
rlabel  s 17 2 17 3 6 C1
port 2 nsew
rlabel  s 17 1 17 2 6 C1
port 2 nsew
rlabel  s 12 22 22 22 6 C1
port 2 nsew
rlabel  s 12 21 22 21 6 C1
port 2 nsew
rlabel  s 12 20 22 20 6 C1
port 2 nsew
rlabel  s 12 18 22 19 6 C1
port 2 nsew
rlabel  s 12 17 22 17 6 C1
port 2 nsew
rlabel  s 12 16 22 16 6 C1
port 2 nsew
rlabel  s 12 14 22 15 6 C1
port 2 nsew
rlabel  s 12 13 22 13 6 C1
port 2 nsew
rlabel  s 12 12 22 12 6 C1
port 2 nsew
rlabel  s 12 11 22 11 6 C1
port 2 nsew
rlabel  s 12 10 22 10 6 C1
port 2 nsew
rlabel  s 12 8 22 9 6 C1
port 2 nsew
rlabel  s 12 7 22 7 6 C1
port 2 nsew
rlabel  s 12 6 22 6 6 C1
port 2 nsew
rlabel  s 12 4 22 5 6 C1
port 2 nsew
rlabel  s 12 3 22 3 6 C1
port 2 nsew
rlabel  s 12 2 22 2 6 C1
port 2 nsew
rlabel  s 12 1 22 1 6 C1
port 2 nsew
rlabel  s 6 21 6 22 6 C1
port 2 nsew
rlabel  s 6 20 6 21 6 C1
port 2 nsew
rlabel  s 6 19 6 20 6 C1
port 2 nsew
rlabel  s 6 17 6 18 6 C1
port 2 nsew
rlabel  s 6 16 6 17 6 C1
port 2 nsew
rlabel  s 6 15 6 16 6 C1
port 2 nsew
rlabel  s 6 13 6 14 6 C1
port 2 nsew
rlabel  s 6 12 6 13 6 C1
port 2 nsew
rlabel  s 6 10 6 11 6 C1
port 2 nsew
rlabel  s 6 9 6 10 6 C1
port 2 nsew
rlabel  s 6 7 6 8 6 C1
port 2 nsew
rlabel  s 6 6 6 7 6 C1
port 2 nsew
rlabel  s 6 5 6 6 6 C1
port 2 nsew
rlabel  s 6 3 6 4 6 C1
port 2 nsew
rlabel  s 6 2 6 3 6 C1
port 2 nsew
rlabel  s 6 1 6 2 6 C1
port 2 nsew
rlabel  s 1 22 11 22 6 C1
port 2 nsew
rlabel  s 1 21 11 21 6 C1
port 2 nsew
rlabel  s 1 20 11 20 6 C1
port 2 nsew
rlabel  s 1 18 11 19 6 C1
port 2 nsew
rlabel  s 1 17 11 17 6 C1
port 2 nsew
rlabel  s 1 16 11 16 6 C1
port 2 nsew
rlabel  s 1 14 11 15 6 C1
port 2 nsew
rlabel  s 1 13 11 13 6 C1
port 2 nsew
rlabel  s 1 12 11 12 6 C1
port 2 nsew
rlabel  s 1 11 11 11 6 C1
port 2 nsew
rlabel  s 1 10 11 10 6 C1
port 2 nsew
rlabel  s 1 8 11 9 6 C1
port 2 nsew
rlabel  s 1 7 11 7 6 C1
port 2 nsew
rlabel  s 1 6 11 6 6 C1
port 2 nsew
rlabel  s 1 4 11 5 6 C1
port 2 nsew
rlabel  s 1 3 11 3 6 C1
port 2 nsew
rlabel  s 1 2 11 2 6 C1
port 2 nsew
rlabel  s 1 1 11 1 6 C1
port 2 nsew
rlabel r s 0 0 22 23 6 M5
port 3 nsew
rlabel metal_blue s 6 6 6 6 6 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22 23
string LEFview TRUE
<< end >>
