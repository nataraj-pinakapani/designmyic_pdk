magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 14 21 1460 203
rect 29 -17 63 21
<< scnmos >>
rect 92 47 122 177
rect 176 47 206 177
rect 260 47 290 177
rect 344 47 374 177
rect 428 47 458 177
rect 512 47 542 177
rect 596 47 626 177
rect 680 47 710 177
rect 764 47 794 177
rect 848 47 878 177
rect 932 47 962 177
rect 1016 47 1046 177
rect 1100 47 1130 177
rect 1184 47 1214 177
rect 1268 47 1298 177
rect 1352 47 1382 177
<< scpmoshvt >>
rect 92 297 122 497
rect 176 297 206 497
rect 260 297 290 497
rect 344 297 374 497
rect 428 297 458 497
rect 512 297 542 497
rect 596 297 626 497
rect 680 297 710 497
rect 764 297 794 497
rect 848 297 878 497
rect 932 297 962 497
rect 1016 297 1046 497
rect 1100 297 1130 497
rect 1184 297 1214 497
rect 1268 297 1298 497
rect 1352 297 1382 497
<< ndiff >>
rect 40 161 92 177
rect 40 127 48 161
rect 82 127 92 161
rect 40 93 92 127
rect 40 59 48 93
rect 82 59 92 93
rect 40 47 92 59
rect 122 161 176 177
rect 122 127 132 161
rect 166 127 176 161
rect 122 93 176 127
rect 122 59 132 93
rect 166 59 176 93
rect 122 47 176 59
rect 206 93 260 177
rect 206 59 216 93
rect 250 59 260 93
rect 206 47 260 59
rect 290 161 344 177
rect 290 127 300 161
rect 334 127 344 161
rect 290 93 344 127
rect 290 59 300 93
rect 334 59 344 93
rect 290 47 344 59
rect 374 93 428 177
rect 374 59 384 93
rect 418 59 428 93
rect 374 47 428 59
rect 458 161 512 177
rect 458 127 468 161
rect 502 127 512 161
rect 458 93 512 127
rect 458 59 468 93
rect 502 59 512 93
rect 458 47 512 59
rect 542 93 596 177
rect 542 59 552 93
rect 586 59 596 93
rect 542 47 596 59
rect 626 161 680 177
rect 626 127 636 161
rect 670 127 680 161
rect 626 93 680 127
rect 626 59 636 93
rect 670 59 680 93
rect 626 47 680 59
rect 710 93 764 177
rect 710 59 720 93
rect 754 59 764 93
rect 710 47 764 59
rect 794 161 848 177
rect 794 127 804 161
rect 838 127 848 161
rect 794 93 848 127
rect 794 59 804 93
rect 838 59 848 93
rect 794 47 848 59
rect 878 93 932 177
rect 878 59 888 93
rect 922 59 932 93
rect 878 47 932 59
rect 962 161 1016 177
rect 962 127 972 161
rect 1006 127 1016 161
rect 962 93 1016 127
rect 962 59 972 93
rect 1006 59 1016 93
rect 962 47 1016 59
rect 1046 93 1100 177
rect 1046 59 1056 93
rect 1090 59 1100 93
rect 1046 47 1100 59
rect 1130 161 1184 177
rect 1130 127 1140 161
rect 1174 127 1184 161
rect 1130 93 1184 127
rect 1130 59 1140 93
rect 1174 59 1184 93
rect 1130 47 1184 59
rect 1214 93 1268 177
rect 1214 59 1224 93
rect 1258 59 1268 93
rect 1214 47 1268 59
rect 1298 161 1352 177
rect 1298 127 1308 161
rect 1342 127 1352 161
rect 1298 93 1352 127
rect 1298 59 1308 93
rect 1342 59 1352 93
rect 1298 47 1352 59
rect 1382 161 1434 177
rect 1382 127 1392 161
rect 1426 127 1434 161
rect 1382 93 1434 127
rect 1382 59 1392 93
rect 1426 59 1434 93
rect 1382 47 1434 59
<< pdiff >>
rect 40 485 92 497
rect 40 451 48 485
rect 82 451 92 485
rect 40 417 92 451
rect 40 383 48 417
rect 82 383 92 417
rect 40 347 92 383
rect 40 313 48 347
rect 82 313 92 347
rect 40 297 92 313
rect 122 485 176 497
rect 122 451 132 485
rect 166 451 176 485
rect 122 417 176 451
rect 122 383 132 417
rect 166 383 176 417
rect 122 347 176 383
rect 122 313 132 347
rect 166 313 176 347
rect 122 297 176 313
rect 206 485 260 497
rect 206 451 216 485
rect 250 451 260 485
rect 206 417 260 451
rect 206 383 216 417
rect 250 383 260 417
rect 206 297 260 383
rect 290 485 344 497
rect 290 451 300 485
rect 334 451 344 485
rect 290 417 344 451
rect 290 383 300 417
rect 334 383 344 417
rect 290 347 344 383
rect 290 313 300 347
rect 334 313 344 347
rect 290 297 344 313
rect 374 485 428 497
rect 374 451 384 485
rect 418 451 428 485
rect 374 417 428 451
rect 374 383 384 417
rect 418 383 428 417
rect 374 297 428 383
rect 458 485 512 497
rect 458 451 468 485
rect 502 451 512 485
rect 458 417 512 451
rect 458 383 468 417
rect 502 383 512 417
rect 458 347 512 383
rect 458 313 468 347
rect 502 313 512 347
rect 458 297 512 313
rect 542 485 596 497
rect 542 451 552 485
rect 586 451 596 485
rect 542 417 596 451
rect 542 383 552 417
rect 586 383 596 417
rect 542 297 596 383
rect 626 485 680 497
rect 626 451 636 485
rect 670 451 680 485
rect 626 417 680 451
rect 626 383 636 417
rect 670 383 680 417
rect 626 347 680 383
rect 626 313 636 347
rect 670 313 680 347
rect 626 297 680 313
rect 710 485 764 497
rect 710 451 720 485
rect 754 451 764 485
rect 710 417 764 451
rect 710 383 720 417
rect 754 383 764 417
rect 710 297 764 383
rect 794 485 848 497
rect 794 451 804 485
rect 838 451 848 485
rect 794 417 848 451
rect 794 383 804 417
rect 838 383 848 417
rect 794 347 848 383
rect 794 313 804 347
rect 838 313 848 347
rect 794 297 848 313
rect 878 485 932 497
rect 878 451 888 485
rect 922 451 932 485
rect 878 417 932 451
rect 878 383 888 417
rect 922 383 932 417
rect 878 297 932 383
rect 962 485 1016 497
rect 962 451 972 485
rect 1006 451 1016 485
rect 962 417 1016 451
rect 962 383 972 417
rect 1006 383 1016 417
rect 962 347 1016 383
rect 962 313 972 347
rect 1006 313 1016 347
rect 962 297 1016 313
rect 1046 485 1100 497
rect 1046 451 1056 485
rect 1090 451 1100 485
rect 1046 417 1100 451
rect 1046 383 1056 417
rect 1090 383 1100 417
rect 1046 297 1100 383
rect 1130 485 1184 497
rect 1130 451 1140 485
rect 1174 451 1184 485
rect 1130 417 1184 451
rect 1130 383 1140 417
rect 1174 383 1184 417
rect 1130 347 1184 383
rect 1130 313 1140 347
rect 1174 313 1184 347
rect 1130 297 1184 313
rect 1214 485 1268 497
rect 1214 451 1224 485
rect 1258 451 1268 485
rect 1214 417 1268 451
rect 1214 383 1224 417
rect 1258 383 1268 417
rect 1214 297 1268 383
rect 1298 485 1352 497
rect 1298 451 1308 485
rect 1342 451 1352 485
rect 1298 417 1352 451
rect 1298 383 1308 417
rect 1342 383 1352 417
rect 1298 347 1352 383
rect 1298 313 1308 347
rect 1342 313 1352 347
rect 1298 297 1352 313
rect 1382 485 1434 497
rect 1382 451 1392 485
rect 1426 451 1434 485
rect 1382 417 1434 451
rect 1382 383 1392 417
rect 1426 383 1434 417
rect 1382 297 1434 383
<< ndiffc >>
rect 48 127 82 161
rect 48 59 82 93
rect 132 127 166 161
rect 132 59 166 93
rect 216 59 250 93
rect 300 127 334 161
rect 300 59 334 93
rect 384 59 418 93
rect 468 127 502 161
rect 468 59 502 93
rect 552 59 586 93
rect 636 127 670 161
rect 636 59 670 93
rect 720 59 754 93
rect 804 127 838 161
rect 804 59 838 93
rect 888 59 922 93
rect 972 127 1006 161
rect 972 59 1006 93
rect 1056 59 1090 93
rect 1140 127 1174 161
rect 1140 59 1174 93
rect 1224 59 1258 93
rect 1308 127 1342 161
rect 1308 59 1342 93
rect 1392 127 1426 161
rect 1392 59 1426 93
<< pdiffc >>
rect 48 451 82 485
rect 48 383 82 417
rect 48 313 82 347
rect 132 451 166 485
rect 132 383 166 417
rect 132 313 166 347
rect 216 451 250 485
rect 216 383 250 417
rect 300 451 334 485
rect 300 383 334 417
rect 300 313 334 347
rect 384 451 418 485
rect 384 383 418 417
rect 468 451 502 485
rect 468 383 502 417
rect 468 313 502 347
rect 552 451 586 485
rect 552 383 586 417
rect 636 451 670 485
rect 636 383 670 417
rect 636 313 670 347
rect 720 451 754 485
rect 720 383 754 417
rect 804 451 838 485
rect 804 383 838 417
rect 804 313 838 347
rect 888 451 922 485
rect 888 383 922 417
rect 972 451 1006 485
rect 972 383 1006 417
rect 972 313 1006 347
rect 1056 451 1090 485
rect 1056 383 1090 417
rect 1140 451 1174 485
rect 1140 383 1174 417
rect 1140 313 1174 347
rect 1224 451 1258 485
rect 1224 383 1258 417
rect 1308 451 1342 485
rect 1308 383 1342 417
rect 1308 313 1342 347
rect 1392 451 1426 485
rect 1392 383 1426 417
<< poly >>
rect 92 497 122 523
rect 176 497 206 523
rect 260 497 290 523
rect 344 497 374 523
rect 428 497 458 523
rect 512 497 542 523
rect 596 497 626 523
rect 680 497 710 523
rect 764 497 794 523
rect 848 497 878 523
rect 932 497 962 523
rect 1016 497 1046 523
rect 1100 497 1130 523
rect 1184 497 1214 523
rect 1268 497 1298 523
rect 1352 497 1382 523
rect 92 265 122 297
rect 176 265 206 297
rect 260 265 290 297
rect 344 265 374 297
rect 428 265 458 297
rect 512 265 542 297
rect 596 265 626 297
rect 680 265 710 297
rect 764 265 794 297
rect 848 265 878 297
rect 932 265 962 297
rect 1016 265 1046 297
rect 1100 265 1130 297
rect 1184 265 1214 297
rect 1268 265 1298 297
rect 1352 265 1382 297
rect 26 249 1382 265
rect 26 215 42 249
rect 76 215 216 249
rect 250 215 384 249
rect 418 215 553 249
rect 587 215 720 249
rect 754 215 888 249
rect 922 215 1055 249
rect 1089 215 1382 249
rect 26 199 1382 215
rect 92 177 122 199
rect 176 177 206 199
rect 260 177 290 199
rect 344 177 374 199
rect 428 177 458 199
rect 512 177 542 199
rect 596 177 626 199
rect 680 177 710 199
rect 764 177 794 199
rect 848 177 878 199
rect 932 177 962 199
rect 1016 177 1046 199
rect 1100 177 1130 199
rect 1184 177 1214 199
rect 1268 177 1298 199
rect 1352 177 1382 199
rect 92 21 122 47
rect 176 21 206 47
rect 260 21 290 47
rect 344 21 374 47
rect 428 21 458 47
rect 512 21 542 47
rect 596 21 626 47
rect 680 21 710 47
rect 764 21 794 47
rect 848 21 878 47
rect 932 21 962 47
rect 1016 21 1046 47
rect 1100 21 1130 47
rect 1184 21 1214 47
rect 1268 21 1298 47
rect 1352 21 1382 47
<< polycont >>
rect 42 215 76 249
rect 216 215 250 249
rect 384 215 418 249
rect 553 215 587 249
rect 720 215 754 249
rect 888 215 922 249
rect 1055 215 1089 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 40 485 82 527
rect 40 451 48 485
rect 40 417 82 451
rect 40 383 48 417
rect 40 347 82 383
rect 40 313 48 347
rect 40 297 82 313
rect 116 485 182 493
rect 116 451 132 485
rect 166 451 182 485
rect 116 417 182 451
rect 116 383 132 417
rect 166 383 182 417
rect 116 347 182 383
rect 216 485 250 527
rect 216 417 250 451
rect 216 367 250 383
rect 284 485 350 493
rect 284 451 300 485
rect 334 451 350 485
rect 284 417 350 451
rect 284 383 300 417
rect 334 383 350 417
rect 116 313 132 347
rect 166 333 182 347
rect 284 347 350 383
rect 384 485 418 527
rect 384 417 418 451
rect 384 367 418 383
rect 452 485 518 493
rect 452 451 468 485
rect 502 451 518 485
rect 452 417 518 451
rect 452 383 468 417
rect 502 383 518 417
rect 284 333 300 347
rect 166 313 300 333
rect 334 333 350 347
rect 452 347 518 383
rect 552 485 586 527
rect 552 417 586 451
rect 552 367 586 383
rect 620 485 686 493
rect 620 451 636 485
rect 670 451 686 485
rect 620 417 686 451
rect 620 383 636 417
rect 670 383 686 417
rect 452 333 468 347
rect 334 313 468 333
rect 502 333 518 347
rect 620 347 686 383
rect 720 485 754 527
rect 720 417 754 451
rect 720 367 754 383
rect 788 485 854 493
rect 788 451 804 485
rect 838 451 854 485
rect 788 417 854 451
rect 788 383 804 417
rect 838 383 854 417
rect 620 333 636 347
rect 502 313 636 333
rect 670 333 686 347
rect 788 347 854 383
rect 888 485 922 527
rect 888 417 922 451
rect 888 367 922 383
rect 956 485 1022 493
rect 956 451 972 485
rect 1006 451 1022 485
rect 956 417 1022 451
rect 956 383 972 417
rect 1006 383 1022 417
rect 788 333 804 347
rect 670 313 804 333
rect 838 333 854 347
rect 956 347 1022 383
rect 1056 485 1090 527
rect 1056 417 1090 451
rect 1056 367 1090 383
rect 1124 485 1190 493
rect 1124 451 1140 485
rect 1174 451 1190 485
rect 1124 417 1190 451
rect 1124 383 1140 417
rect 1174 383 1190 417
rect 956 333 972 347
rect 838 313 972 333
rect 1006 333 1022 347
rect 1124 347 1190 383
rect 1224 485 1258 527
rect 1224 417 1258 451
rect 1224 367 1258 383
rect 1292 485 1358 493
rect 1292 451 1308 485
rect 1342 451 1358 485
rect 1292 417 1358 451
rect 1292 383 1308 417
rect 1342 383 1358 417
rect 1124 333 1140 347
rect 1006 313 1140 333
rect 1174 333 1190 347
rect 1292 347 1358 383
rect 1392 485 1434 527
rect 1426 451 1434 485
rect 1392 417 1434 451
rect 1426 383 1434 417
rect 1392 367 1434 383
rect 1292 333 1308 347
rect 1174 313 1308 333
rect 1342 313 1358 347
rect 116 299 1358 313
rect 17 249 1105 263
rect 17 215 42 249
rect 76 215 216 249
rect 250 215 384 249
rect 418 215 553 249
rect 587 215 720 249
rect 754 215 888 249
rect 922 215 1055 249
rect 1089 215 1105 249
rect 1292 181 1358 299
rect 36 161 82 177
rect 36 127 48 161
rect 36 93 82 127
rect 36 59 48 93
rect 36 17 82 59
rect 116 161 1358 181
rect 116 127 132 161
rect 166 143 300 161
rect 166 127 182 143
rect 116 93 182 127
rect 284 127 300 143
rect 334 143 468 161
rect 334 127 350 143
rect 116 59 132 93
rect 166 59 182 93
rect 116 51 182 59
rect 216 93 250 109
rect 216 17 250 59
rect 284 93 350 127
rect 452 127 468 143
rect 502 143 636 161
rect 502 127 518 143
rect 284 59 300 93
rect 334 59 350 93
rect 284 51 350 59
rect 384 93 418 109
rect 384 17 418 59
rect 452 93 518 127
rect 620 127 636 143
rect 670 143 804 161
rect 670 127 686 143
rect 452 59 468 93
rect 502 59 518 93
rect 452 51 518 59
rect 552 93 586 109
rect 552 17 586 59
rect 620 93 686 127
rect 788 127 804 143
rect 838 143 972 161
rect 838 127 854 143
rect 620 59 636 93
rect 670 59 686 93
rect 620 51 686 59
rect 720 93 754 109
rect 720 17 754 59
rect 788 93 854 127
rect 956 127 972 143
rect 1006 143 1140 161
rect 1006 127 1022 143
rect 788 59 804 93
rect 838 59 854 93
rect 788 51 854 59
rect 888 93 922 109
rect 888 17 922 59
rect 956 93 1022 127
rect 1124 127 1140 143
rect 1174 143 1308 161
rect 1174 127 1190 143
rect 956 59 972 93
rect 1006 59 1022 93
rect 956 51 1022 59
rect 1056 93 1090 109
rect 1056 17 1090 59
rect 1124 93 1190 127
rect 1292 127 1308 143
rect 1342 127 1358 161
rect 1124 59 1140 93
rect 1174 59 1190 93
rect 1124 51 1190 59
rect 1224 93 1258 109
rect 1224 17 1258 59
rect 1292 93 1358 127
rect 1292 59 1308 93
rect 1342 59 1358 93
rect 1292 51 1358 59
rect 1392 161 1434 177
rect 1426 127 1434 161
rect 1392 93 1434 127
rect 1426 59 1434 93
rect 1392 17 1434 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 1317 221 1351 255 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 1317 153 1351 187 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 inv_16
rlabel metal1 s 0 -48 1472 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 2246974
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 2235486
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 36.800 0.000 
<< end >>
