magic
tech minimum
timestamp 1644097874
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -4 -4 4 19
string LEFview TRUE
<< end >>
