/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/fixed_devices/sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18_fail.cdl