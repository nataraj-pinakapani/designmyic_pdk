magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 16 21 1159 203
rect 29 -17 63 21
<< locali >>
rect 121 257 177 341
rect 85 215 177 257
rect 211 289 445 341
rect 211 181 291 289
rect 211 145 445 181
rect 756 215 964 255
rect 998 215 1179 255
rect 211 51 277 145
rect 379 51 445 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 409 87 493
rect 127 443 193 527
rect 295 443 361 527
rect 463 443 529 527
rect 17 375 513 409
rect 17 291 87 375
rect 17 171 51 291
rect 479 323 513 375
rect 563 393 597 493
rect 640 427 690 527
rect 737 459 953 493
rect 737 427 785 459
rect 827 393 876 425
rect 563 359 876 393
rect 479 289 581 323
rect 325 215 513 255
rect 547 249 581 289
rect 547 215 627 249
rect 17 53 109 171
rect 143 17 177 181
rect 479 179 513 215
rect 679 179 717 359
rect 827 289 876 359
rect 919 333 953 459
rect 987 367 1053 527
rect 1087 333 1142 493
rect 919 291 1142 333
rect 479 145 717 179
rect 311 17 345 111
rect 647 129 717 145
rect 751 145 1142 181
rect 479 17 513 111
rect 751 95 801 145
rect 561 51 801 95
rect 835 17 869 111
rect 903 51 969 145
rect 1003 17 1037 111
rect 1071 53 1142 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 998 215 1179 255 6 A1
port 1 nsew signal input
rlabel locali s 756 215 964 255 6 A2
port 2 nsew signal input
rlabel locali s 85 215 177 257 6 B1_N
port 3 nsew signal input
rlabel locali s 121 257 177 341 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 16 21 1159 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 379 51 445 145 6 X
port 8 nsew signal output
rlabel locali s 211 51 277 145 6 X
port 8 nsew signal output
rlabel locali s 211 145 445 181 6 X
port 8 nsew signal output
rlabel locali s 211 181 291 289 6 X
port 8 nsew signal output
rlabel locali s 211 289 445 341 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1328502
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1319502
<< end >>
