magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< locali >>
rect 0 792 788 826
rect 822 797 876 826
rect 0 772 54 792
rect 0 738 10 772
rect 44 738 54 772
rect 822 763 832 797
rect 866 763 876 797
rect 822 756 876 763
rect 0 700 54 738
rect 88 725 876 756
rect 88 722 832 725
rect 0 666 10 700
rect 44 686 54 700
rect 822 691 832 722
rect 866 691 876 725
rect 44 666 788 686
rect 0 652 788 666
rect 822 653 876 691
rect 0 628 54 652
rect 0 594 10 628
rect 44 594 54 628
rect 822 619 832 653
rect 866 619 876 653
rect 822 616 876 619
rect 0 556 54 594
rect 88 582 876 616
rect 0 522 10 556
rect 44 546 54 556
rect 822 581 876 582
rect 822 547 832 581
rect 866 547 876 581
rect 44 522 788 546
rect 0 512 788 522
rect 0 484 54 512
rect 0 450 10 484
rect 44 450 54 484
rect 822 509 876 547
rect 822 476 832 509
rect 0 412 54 450
rect 88 475 832 476
rect 866 475 876 509
rect 88 442 876 475
rect 0 378 10 412
rect 44 406 54 412
rect 822 437 876 442
rect 44 378 788 406
rect 0 372 788 378
rect 822 403 832 437
rect 866 403 876 437
rect 0 340 54 372
rect 0 306 10 340
rect 44 306 54 340
rect 822 365 876 403
rect 822 336 832 365
rect 0 268 54 306
rect 88 331 832 336
rect 866 331 876 365
rect 88 302 876 331
rect 0 234 10 268
rect 44 266 54 268
rect 822 293 876 302
rect 44 234 788 266
rect 0 232 788 234
rect 822 259 832 293
rect 866 259 876 293
rect 0 196 54 232
rect 822 221 876 259
rect 822 196 832 221
rect 0 162 10 196
rect 44 162 54 196
rect 88 187 832 196
rect 866 187 876 221
rect 88 162 876 187
rect 0 126 54 162
rect 822 149 876 162
rect 0 124 788 126
rect 0 90 10 124
rect 44 92 788 124
rect 822 115 832 149
rect 866 115 876 149
rect 822 92 876 115
rect 44 90 54 92
rect 0 64 54 90
<< viali >>
rect 10 738 44 772
rect 832 763 866 797
rect 10 666 44 700
rect 832 691 866 725
rect 10 594 44 628
rect 832 619 866 653
rect 10 522 44 556
rect 832 547 866 581
rect 10 450 44 484
rect 832 475 866 509
rect 10 378 44 412
rect 832 403 866 437
rect 10 306 44 340
rect 832 331 866 365
rect 10 234 44 268
rect 832 259 866 293
rect 10 162 44 196
rect 832 187 866 221
rect 10 90 44 124
rect 832 115 866 149
<< metal1 >>
rect 0 912 876 918
rect 0 860 76 912
rect 128 860 140 912
rect 192 860 204 912
rect 256 860 268 912
rect 320 860 332 912
rect 384 860 396 912
rect 448 860 460 912
rect 512 860 524 912
rect 576 860 588 912
rect 640 860 652 912
rect 704 860 716 912
rect 768 860 876 912
rect 0 854 876 860
rect 0 809 54 826
rect 0 757 1 809
rect 53 757 54 809
rect 0 745 10 757
rect 44 745 54 757
rect 0 693 1 745
rect 53 693 54 745
rect 0 681 10 693
rect 44 681 54 693
rect 0 629 1 681
rect 53 629 54 681
rect 0 628 54 629
rect 0 617 10 628
rect 44 617 54 628
rect 0 565 1 617
rect 53 565 54 617
rect 0 556 54 565
rect 0 553 10 556
rect 44 553 54 556
rect 0 501 1 553
rect 53 501 54 553
rect 0 489 54 501
rect 0 437 1 489
rect 53 437 54 489
rect 0 425 54 437
rect 0 373 1 425
rect 53 373 54 425
rect 0 361 54 373
rect 0 309 1 361
rect 53 309 54 361
rect 0 306 10 309
rect 44 306 54 309
rect 0 297 54 306
rect 0 245 1 297
rect 53 245 54 297
rect 0 234 10 245
rect 44 234 54 245
rect 0 233 54 234
rect 0 181 1 233
rect 53 181 54 233
rect 0 169 10 181
rect 44 169 54 181
rect 0 117 1 169
rect 53 117 54 169
rect 0 105 10 117
rect 44 105 54 117
rect 0 53 1 105
rect 53 64 54 105
rect 88 64 116 826
rect 144 92 172 854
rect 200 64 228 826
rect 256 92 284 854
rect 312 64 340 826
rect 368 92 396 854
rect 424 64 452 826
rect 480 92 508 854
rect 536 64 564 826
rect 592 92 620 854
rect 648 64 676 826
rect 704 92 732 854
rect 760 64 788 826
rect 822 797 876 854
rect 822 790 832 797
rect 866 790 876 797
rect 822 738 823 790
rect 875 738 876 790
rect 822 726 876 738
rect 822 674 823 726
rect 875 674 876 726
rect 822 662 876 674
rect 822 610 823 662
rect 875 610 876 662
rect 822 598 876 610
rect 822 546 823 598
rect 875 546 876 598
rect 822 534 876 546
rect 822 482 823 534
rect 875 482 876 534
rect 822 475 832 482
rect 866 475 876 482
rect 822 470 876 475
rect 822 418 823 470
rect 875 418 876 470
rect 822 406 832 418
rect 866 406 876 418
rect 822 354 823 406
rect 875 354 876 406
rect 822 342 832 354
rect 866 342 876 354
rect 822 290 823 342
rect 875 290 876 342
rect 822 278 832 290
rect 866 278 876 290
rect 822 226 823 278
rect 875 226 876 278
rect 822 221 876 226
rect 822 214 832 221
rect 866 214 876 221
rect 822 162 823 214
rect 875 162 876 214
rect 822 150 876 162
rect 822 98 823 150
rect 875 98 876 150
rect 822 92 876 98
rect 53 58 876 64
rect 53 53 76 58
rect 0 6 76 53
rect 128 6 140 58
rect 192 6 204 58
rect 256 6 268 58
rect 320 6 332 58
rect 384 6 396 58
rect 448 6 460 58
rect 512 6 524 58
rect 576 6 588 58
rect 640 6 652 58
rect 704 6 716 58
rect 768 6 876 58
rect 0 0 876 6
<< via1 >>
rect 76 860 128 912
rect 140 860 192 912
rect 204 860 256 912
rect 268 860 320 912
rect 332 860 384 912
rect 396 860 448 912
rect 460 860 512 912
rect 524 860 576 912
rect 588 860 640 912
rect 652 860 704 912
rect 716 860 768 912
rect 1 772 53 809
rect 1 757 10 772
rect 10 757 44 772
rect 44 757 53 772
rect 1 738 10 745
rect 10 738 44 745
rect 44 738 53 745
rect 1 700 53 738
rect 1 693 10 700
rect 10 693 44 700
rect 44 693 53 700
rect 1 666 10 681
rect 10 666 44 681
rect 44 666 53 681
rect 1 629 53 666
rect 1 594 10 617
rect 10 594 44 617
rect 44 594 53 617
rect 1 565 53 594
rect 1 522 10 553
rect 10 522 44 553
rect 44 522 53 553
rect 1 501 53 522
rect 1 484 53 489
rect 1 450 10 484
rect 10 450 44 484
rect 44 450 53 484
rect 1 437 53 450
rect 1 412 53 425
rect 1 378 10 412
rect 10 378 44 412
rect 44 378 53 412
rect 1 373 53 378
rect 1 340 53 361
rect 1 309 10 340
rect 10 309 44 340
rect 44 309 53 340
rect 1 268 53 297
rect 1 245 10 268
rect 10 245 44 268
rect 44 245 53 268
rect 1 196 53 233
rect 1 181 10 196
rect 10 181 44 196
rect 44 181 53 196
rect 1 162 10 169
rect 10 162 44 169
rect 44 162 53 169
rect 1 124 53 162
rect 1 117 10 124
rect 10 117 44 124
rect 44 117 53 124
rect 1 90 10 105
rect 10 90 44 105
rect 44 90 53 105
rect 1 53 53 90
rect 823 763 832 790
rect 832 763 866 790
rect 866 763 875 790
rect 823 738 875 763
rect 823 725 875 726
rect 823 691 832 725
rect 832 691 866 725
rect 866 691 875 725
rect 823 674 875 691
rect 823 653 875 662
rect 823 619 832 653
rect 832 619 866 653
rect 866 619 875 653
rect 823 610 875 619
rect 823 581 875 598
rect 823 547 832 581
rect 832 547 866 581
rect 866 547 875 581
rect 823 546 875 547
rect 823 509 875 534
rect 823 482 832 509
rect 832 482 866 509
rect 866 482 875 509
rect 823 437 875 470
rect 823 418 832 437
rect 832 418 866 437
rect 866 418 875 437
rect 823 403 832 406
rect 832 403 866 406
rect 866 403 875 406
rect 823 365 875 403
rect 823 354 832 365
rect 832 354 866 365
rect 866 354 875 365
rect 823 331 832 342
rect 832 331 866 342
rect 866 331 875 342
rect 823 293 875 331
rect 823 290 832 293
rect 832 290 866 293
rect 866 290 875 293
rect 823 259 832 278
rect 832 259 866 278
rect 866 259 875 278
rect 823 226 875 259
rect 823 187 832 214
rect 832 187 866 214
rect 866 187 875 214
rect 823 162 875 187
rect 823 149 875 150
rect 823 115 832 149
rect 832 115 866 149
rect 866 115 875 149
rect 823 98 875 115
rect 76 6 128 58
rect 140 6 192 58
rect 204 6 256 58
rect 268 6 320 58
rect 332 6 384 58
rect 396 6 448 58
rect 460 6 512 58
rect 524 6 576 58
rect 588 6 640 58
rect 652 6 704 58
rect 716 6 768 58
<< metal2 >>
rect 0 912 876 918
rect 0 860 76 912
rect 128 860 140 912
rect 192 860 204 912
rect 256 860 268 912
rect 320 860 332 912
rect 384 860 396 912
rect 448 860 460 912
rect 512 860 524 912
rect 576 860 588 912
rect 640 860 652 912
rect 704 860 716 912
rect 768 860 876 912
rect 0 854 876 860
rect 0 809 54 826
rect 0 757 1 809
rect 53 757 54 809
rect 0 745 54 757
rect 0 693 1 745
rect 53 693 54 745
rect 0 681 54 693
rect 0 629 1 681
rect 53 629 54 681
rect 0 617 54 629
rect 0 565 1 617
rect 53 565 54 617
rect 0 553 54 565
rect 0 501 1 553
rect 53 501 54 553
rect 0 489 54 501
rect 0 437 1 489
rect 53 437 54 489
rect 0 425 54 437
rect 0 373 1 425
rect 53 373 54 425
rect 0 361 54 373
rect 0 309 1 361
rect 53 309 54 361
rect 0 297 54 309
rect 0 245 1 297
rect 53 245 54 297
rect 0 233 54 245
rect 0 181 1 233
rect 53 181 54 233
rect 0 169 54 181
rect 0 117 1 169
rect 53 117 54 169
rect 0 105 54 117
rect 0 53 1 105
rect 53 64 54 105
rect 88 92 116 854
rect 144 64 172 826
rect 200 92 228 854
rect 256 64 284 826
rect 312 92 340 854
rect 368 64 396 826
rect 424 92 452 854
rect 480 64 508 826
rect 536 92 564 854
rect 592 64 620 826
rect 648 92 676 854
rect 704 64 732 826
rect 760 92 788 854
rect 822 790 876 854
rect 822 738 823 790
rect 875 738 876 790
rect 822 726 876 738
rect 822 674 823 726
rect 875 674 876 726
rect 822 662 876 674
rect 822 610 823 662
rect 875 610 876 662
rect 822 598 876 610
rect 822 546 823 598
rect 875 546 876 598
rect 822 534 876 546
rect 822 482 823 534
rect 875 482 876 534
rect 822 470 876 482
rect 822 418 823 470
rect 875 418 876 470
rect 822 406 876 418
rect 822 354 823 406
rect 875 354 876 406
rect 822 342 876 354
rect 822 290 823 342
rect 875 290 876 342
rect 822 278 876 290
rect 822 226 823 278
rect 875 226 876 278
rect 822 214 876 226
rect 822 162 823 214
rect 875 162 876 214
rect 822 150 876 162
rect 822 98 823 150
rect 875 98 876 150
rect 822 92 876 98
rect 53 58 876 64
rect 53 53 76 58
rect 0 6 76 53
rect 128 6 140 58
rect 192 6 204 58
rect 256 6 268 58
rect 320 6 332 58
rect 384 6 396 58
rect 448 6 460 58
rect 512 6 524 58
rect 576 6 588 58
rect 640 6 652 58
rect 704 6 716 58
rect 768 6 876 58
rect 0 0 876 6
<< labels >>
flabel comment s 807 460 807 460 0 FreeSans 200 180 0 0 B
flabel comment s 807 180 807 180 0 FreeSans 200 180 0 0 B
flabel comment s 807 320 807 320 0 FreeSans 200 180 0 0 B
flabel comment s 807 740 807 740 0 FreeSans 200 180 0 0 B
flabel comment s 807 600 807 600 0 FreeSans 200 180 0 0 B
flabel comment s 63 670 63 670 0 FreeSans 200 0 0 0 A
flabel comment s 63 250 63 250 0 FreeSans 200 0 0 0 A
flabel comment s 63 810 63 810 0 FreeSans 200 0 0 0 A
flabel comment s 63 110 63 110 0 FreeSans 200 0 0 0 A
flabel comment s 63 390 63 390 0 FreeSans 200 0 0 0 A
flabel comment s 63 530 63 530 0 FreeSans 200 0 0 0 A
flabel comment s 103 839 103 839 0 FreeSans 200 0 0 0 B
flabel comment s 215 839 215 839 0 FreeSans 200 0 0 0 B
flabel comment s 327 839 327 839 0 FreeSans 200 0 0 0 B
flabel comment s 439 839 439 839 0 FreeSans 200 0 0 0 B
flabel comment s 551 839 551 839 0 FreeSans 200 0 0 0 B
flabel comment s 663 839 663 839 0 FreeSans 200 0 0 0 B
flabel comment s 775 839 775 839 0 FreeSans 200 0 0 0 B
flabel comment s 719 79 719 79 0 FreeSans 200 0 0 0 A
flabel comment s 156 839 156 839 0 FreeSans 200 0 0 0 B
flabel comment s 268 839 268 839 0 FreeSans 200 0 0 0 B
flabel comment s 380 839 380 839 0 FreeSans 200 0 0 0 B
flabel comment s 492 839 492 839 0 FreeSans 200 0 0 0 B
flabel comment s 604 839 604 839 0 FreeSans 200 0 0 0 B
flabel comment s 716 839 716 839 0 FreeSans 200 0 0 0 B
flabel comment s 103 79 103 79 0 FreeSans 200 0 0 0 A
flabel comment s 215 79 215 79 0 FreeSans 200 0 0 0 A
flabel comment s 327 79 327 79 0 FreeSans 200 0 0 0 A
flabel comment s 439 79 439 79 0 FreeSans 200 0 0 0 A
flabel comment s 551 79 551 79 0 FreeSans 200 0 0 0 A
flabel comment s 663 79 663 79 0 FreeSans 200 0 0 0 A
flabel comment s 775 79 775 79 0 FreeSans 200 0 0 0 A
flabel comment s 495 79 495 79 0 FreeSans 200 0 0 0 A
flabel comment s 607 79 607 79 0 FreeSans 200 0 0 0 A
flabel comment s 159 79 159 79 0 FreeSans 200 0 0 0 A
flabel comment s 271 79 271 79 0 FreeSans 200 0 0 0 A
flabel comment s 383 79 383 79 0 FreeSans 200 0 0 0 A
<< properties >>
string GDS_END 70294
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 60000
<< end >>
