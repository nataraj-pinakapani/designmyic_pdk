/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__rf_pfet_01v8_aF02W2p00L0p15.spice