/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_e/begin_of_life/mm.spice