magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< obsli1 >>
rect 0 2272 4498 2338
rect 0 66 28 2244
rect 56 94 84 2272
rect 112 66 140 2244
rect 168 94 196 2272
rect 224 66 252 2244
rect 280 94 308 2272
rect 336 66 364 2244
rect 392 94 420 2272
rect 448 66 476 2244
rect 504 94 532 2272
rect 560 66 588 2244
rect 616 94 644 2272
rect 672 66 700 2244
rect 728 94 756 2272
rect 784 66 812 2244
rect 840 94 868 2272
rect 896 66 924 2244
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 1064 94 1092 2272
rect 1120 66 1148 2244
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1288 94 1316 2272
rect 1344 66 1372 2244
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1512 94 1540 2272
rect 1568 66 1596 2244
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1736 94 1764 2272
rect 1792 66 1820 2244
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1960 94 1988 2272
rect 2016 66 2044 2244
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2184 94 2212 2272
rect 2240 66 2268 2244
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2408 94 2436 2272
rect 2464 66 2492 2244
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2632 94 2660 2272
rect 2688 66 2716 2244
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2856 94 2884 2272
rect 2912 66 2940 2244
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 3080 94 3108 2272
rect 3136 66 3164 2244
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3304 94 3332 2272
rect 3360 66 3388 2244
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3528 94 3556 2272
rect 3584 66 3612 2244
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3752 94 3780 2272
rect 3808 66 3836 2244
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3976 94 4004 2272
rect 4032 66 4060 2244
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4200 94 4228 2272
rect 4256 66 4284 2244
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4424 94 4498 2272
rect 0 0 4498 66
<< obsm1 >>
rect 0 2272 4498 2338
rect 0 94 28 2272
rect 56 66 84 2244
rect 112 94 140 2272
rect 168 66 196 2244
rect 224 94 252 2272
rect 280 66 308 2244
rect 336 94 364 2272
rect 392 66 420 2244
rect 448 94 476 2272
rect 504 66 532 2244
rect 560 94 588 2272
rect 616 66 644 2244
rect 672 94 700 2272
rect 728 66 756 2244
rect 784 94 812 2272
rect 840 66 868 2244
rect 896 94 924 2272
rect 952 66 980 2244
rect 1008 94 1036 2272
rect 1064 66 1092 2244
rect 1120 94 1148 2272
rect 1176 66 1204 2244
rect 1232 94 1260 2272
rect 1288 66 1316 2244
rect 1344 94 1372 2272
rect 1400 66 1428 2244
rect 1456 94 1484 2272
rect 1512 66 1540 2244
rect 1568 94 1596 2272
rect 1624 66 1652 2244
rect 1680 94 1708 2272
rect 1736 66 1764 2244
rect 1792 94 1820 2272
rect 1848 66 1876 2244
rect 1904 94 1932 2272
rect 1960 66 1988 2244
rect 2016 94 2044 2272
rect 2072 66 2100 2244
rect 2128 94 2156 2272
rect 2184 66 2212 2244
rect 2240 94 2268 2272
rect 2296 66 2324 2244
rect 2352 94 2380 2272
rect 2408 66 2436 2244
rect 2464 94 2492 2272
rect 2520 66 2548 2244
rect 2576 94 2604 2272
rect 2632 66 2660 2244
rect 2688 94 2716 2272
rect 2744 66 2772 2244
rect 2800 94 2828 2272
rect 2856 66 2884 2244
rect 2912 94 2940 2272
rect 2968 66 2996 2244
rect 3024 94 3052 2272
rect 3080 66 3108 2244
rect 3136 94 3164 2272
rect 3192 66 3220 2244
rect 3248 94 3276 2272
rect 3304 66 3332 2244
rect 3360 94 3388 2272
rect 3416 66 3444 2244
rect 3472 94 3500 2272
rect 3528 66 3556 2244
rect 3584 94 3612 2272
rect 3640 66 3668 2244
rect 3696 94 3724 2272
rect 3752 66 3780 2244
rect 3808 94 3836 2272
rect 3864 66 3892 2244
rect 3920 94 3948 2272
rect 3976 66 4004 2244
rect 4032 94 4060 2272
rect 4088 66 4116 2244
rect 4144 94 4172 2272
rect 4200 66 4228 2244
rect 4256 94 4284 2272
rect 4312 66 4340 2244
rect 4368 94 4396 2272
rect 4424 66 4498 2244
rect 0 0 4498 66
<< obsm2 >>
rect 0 66 28 2338
rect 56 2272 196 2338
rect 56 94 84 2272
rect 112 66 140 2244
rect 0 0 140 66
rect 168 0 196 2272
rect 224 66 252 2338
rect 280 2272 420 2338
rect 280 94 308 2272
rect 336 66 364 2244
rect 224 0 364 66
rect 392 0 420 2272
rect 448 66 476 2338
rect 504 2272 644 2338
rect 504 94 532 2272
rect 560 66 588 2244
rect 448 0 588 66
rect 616 0 644 2272
rect 672 66 700 2338
rect 728 2272 868 2338
rect 728 94 756 2272
rect 784 66 812 2244
rect 672 0 812 66
rect 840 0 868 2272
rect 896 66 924 2338
rect 952 2272 1092 2338
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 896 0 1036 66
rect 1064 0 1092 2272
rect 1120 66 1148 2338
rect 1176 2272 1316 2338
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1120 0 1260 66
rect 1288 0 1316 2272
rect 1344 66 1372 2338
rect 1400 2272 1540 2338
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1344 0 1484 66
rect 1512 0 1540 2272
rect 1568 66 1596 2338
rect 1624 2272 1764 2338
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1568 0 1708 66
rect 1736 0 1764 2272
rect 1792 66 1820 2338
rect 1848 2272 1988 2338
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1792 0 1932 66
rect 1960 0 1988 2272
rect 2016 66 2044 2338
rect 2072 2272 2212 2338
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2016 0 2156 66
rect 2184 0 2212 2272
rect 2240 66 2268 2338
rect 2296 2272 2436 2338
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2240 0 2380 66
rect 2408 0 2436 2272
rect 2464 66 2492 2338
rect 2520 2272 2660 2338
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2464 0 2604 66
rect 2632 0 2660 2272
rect 2688 66 2716 2338
rect 2744 2272 2884 2338
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2688 0 2828 66
rect 2856 0 2884 2272
rect 2912 66 2940 2338
rect 2968 2272 3108 2338
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 2912 0 3052 66
rect 3080 0 3108 2272
rect 3136 66 3164 2338
rect 3192 2272 3332 2338
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3136 0 3276 66
rect 3304 0 3332 2272
rect 3360 66 3388 2338
rect 3416 2272 3556 2338
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3360 0 3500 66
rect 3528 0 3556 2272
rect 3584 66 3612 2338
rect 3640 2272 3780 2338
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3584 0 3724 66
rect 3752 0 3780 2272
rect 3808 66 3836 2338
rect 3864 2272 4004 2338
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3808 0 3948 66
rect 3976 0 4004 2272
rect 4032 66 4060 2338
rect 4088 2272 4498 2338
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4032 0 4172 66
rect 4200 0 4228 2272
rect 4256 66 4284 2244
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4424 94 4498 2272
rect 4256 0 4498 66
<< obsm3 >>
rect 0 2272 4498 2338
rect 0 126 60 2272
rect 120 66 180 2212
rect 240 126 300 2272
rect 360 66 420 2212
rect 480 126 540 2272
rect 600 66 660 2212
rect 720 126 780 2272
rect 840 66 900 2212
rect 960 126 1020 2272
rect 1080 66 1140 2212
rect 1200 126 1260 2272
rect 1320 66 1380 2212
rect 1440 126 1500 2272
rect 1560 66 1620 2212
rect 1680 126 1740 2272
rect 1800 66 1860 2212
rect 1920 126 1980 2272
rect 2040 66 2100 2212
rect 2160 126 2220 2272
rect 2280 66 2340 2212
rect 2400 126 2460 2272
rect 2520 66 2580 2212
rect 2640 126 2700 2272
rect 2760 66 2820 2212
rect 2880 126 2940 2272
rect 3000 66 3060 2212
rect 3120 126 3180 2272
rect 3240 66 3300 2212
rect 3360 126 3420 2272
rect 3480 66 3540 2212
rect 3600 126 3660 2272
rect 3720 66 3780 2212
rect 3840 126 3900 2272
rect 3960 66 4020 2212
rect 4080 126 4140 2272
rect 4200 66 4260 2212
rect 4320 126 4498 2272
rect 0 0 4498 66
<< obsm4 >>
rect 0 2272 4498 2338
rect 0 66 60 2212
rect 120 2027 420 2272
rect 120 126 180 2027
rect 240 311 300 1967
rect 360 371 420 2027
rect 480 311 540 2212
rect 240 66 540 311
rect 600 126 660 2272
rect 720 66 780 2212
rect 840 126 900 2272
rect 960 66 1020 2212
rect 1080 126 1140 2272
rect 1200 66 1260 2212
rect 1320 126 1380 2272
rect 1440 66 1500 2212
rect 1560 2027 1860 2272
rect 1560 126 1620 2027
rect 1680 311 1740 1967
rect 1800 371 1860 2027
rect 1920 311 1980 2212
rect 1680 66 1980 311
rect 2040 126 2100 2272
rect 2160 66 2220 2212
rect 2280 126 2340 2272
rect 2400 66 2460 2212
rect 2520 126 2580 2272
rect 2640 66 2700 2212
rect 2760 126 2820 2272
rect 2880 66 2940 2212
rect 3000 2027 3300 2272
rect 3000 126 3060 2027
rect 3120 311 3180 1967
rect 3240 371 3300 2027
rect 3360 311 3420 2212
rect 3120 66 3420 311
rect 3480 126 3540 2272
rect 3600 66 3660 2212
rect 3720 126 3780 2272
rect 3840 66 3900 2212
rect 3960 126 4020 2272
rect 4080 66 4140 2212
rect 4200 126 4260 2272
rect 4320 66 4498 2212
rect 0 0 4498 66
<< obsm5 >>
rect 0 2003 4498 2338
rect 0 655 320 2003
rect 640 335 960 1683
rect 1280 655 1600 2003
rect 1920 335 2240 1683
rect 2560 655 2880 2003
rect 3200 335 3520 1683
rect 3840 655 4498 2003
rect 0 0 4498 335
<< properties >>
string FIXED_BBOX 0 0 4498 2338
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1495724
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 1432936
<< end >>
