magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 1 0 3 1 8 DRAIN
port 1 nsew
rlabel  s 1 1 3 1 6 GATE
port 2 nsew
rlabel  s 3 0 3 1 8 SOURCE
port 3 nsew
rlabel  s 2 0 2 1 8 SOURCE
port 3 nsew
rlabel  s 1 0 1 1 8 SOURCE
port 3 nsew
rlabel  s 0 0 0 1 2 SOURCE
port 3 nsew
rlabel  s 0 0 3 0 8 SOURCE
port 3 nsew
rlabel metal_blue s 0 1 0 1 4 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 3 2
string LEFview TRUE
<< end >>
