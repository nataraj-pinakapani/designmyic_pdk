magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel 
 s 1 35 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 1 50 24 51 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 51 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 51 50 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 35 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 50 24 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 51 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 51 50 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 46 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 54 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 51 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 50 75 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 50 75 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 38 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 75 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 75 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 36 75 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 36 75 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 35 75 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 35 75 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 51 74 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 50 74 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 50 74 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 38 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 36 74 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 36 74 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 35 74 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 35 74 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 51 74 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 50 74 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 50 74 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 38 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 37 74 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 36 74 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 36 74 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 35 74 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 74 35 74 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 51 73 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 50 73 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 50 73 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 36 73 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 36 73 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 35 73 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 35 73 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 51 73 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 50 73 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 50 73 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 36 73 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 36 73 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 35 73 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 73 35 73 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 51 73 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 50 73 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 50 73 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 73 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 73 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 36 73 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 36 73 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 35 73 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 35 73 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 51 72 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 50 72 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 50 72 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 36 72 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 36 72 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 35 72 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 35 72 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 51 72 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 50 72 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 50 72 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 38 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 37 72 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 36 72 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 36 72 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 35 72 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 72 35 72 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 51 71 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 50 71 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 50 71 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 36 71 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 36 71 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 35 71 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 35 71 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 51 71 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 50 71 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 50 71 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 36 71 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 36 71 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 35 71 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 71 35 71 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 51 71 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 50 71 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 50 71 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 71 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 71 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 36 71 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 36 71 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 35 71 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 35 71 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 51 70 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 50 70 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 50 70 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 36 70 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 36 70 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 35 70 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 35 70 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 51 70 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 50 70 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 50 70 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 38 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 37 70 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 36 70 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 36 70 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 35 70 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 70 35 70 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 51 69 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 50 69 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 50 69 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 36 69 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 36 69 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 35 69 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 35 69 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 51 69 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 50 69 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 50 69 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 38 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 37 69 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 36 69 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 36 69 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 35 69 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 69 35 69 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 51 68 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 50 68 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 50 68 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 36 68 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 36 68 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 35 68 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 35 68 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 51 68 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 50 68 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 50 68 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 38 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 36 68 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 36 68 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 35 68 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 68 35 68 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 51 68 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 50 68 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 50 68 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 38 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 68 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 68 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 36 68 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 36 68 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 35 68 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 35 68 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 51 67 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 50 67 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 50 67 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 36 67 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 36 67 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 35 67 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 35 67 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 51 67 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 50 67 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 50 67 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 38 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 37 67 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 36 67 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 36 67 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 35 67 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 67 35 67 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 51 66 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 50 66 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 50 66 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 38 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 36 66 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 36 66 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 35 66 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 35 66 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 51 66 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 50 66 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 50 66 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 38 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 36 66 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 36 66 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 35 66 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 66 35 66 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 51 66 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 50 66 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 50 66 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 66 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 66 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 36 66 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 36 66 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 35 66 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 35 66 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 51 65 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 50 65 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 50 65 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 36 65 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 36 65 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 35 65 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 35 65 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 51 65 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 50 65 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 50 65 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 38 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 37 65 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 36 65 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 36 65 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 35 65 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 65 35 65 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 51 64 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 50 64 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 50 64 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 36 64 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 36 64 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 35 64 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 35 64 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 51 64 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 50 64 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 50 64 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 36 64 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 36 64 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 35 64 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 64 35 64 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 51 64 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 50 64 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 50 64 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 64 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 64 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 36 64 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 36 64 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 35 64 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 35 64 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 51 63 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 50 63 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 50 63 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 36 63 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 36 63 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 35 63 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 35 63 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 51 63 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 50 63 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 50 63 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 38 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 37 63 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 36 63 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 36 63 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 35 63 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 63 35 63 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 51 62 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 50 62 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 50 62 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 36 62 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 36 62 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 35 62 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 35 62 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 51 62 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 50 62 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 50 62 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 36 62 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 36 62 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 35 62 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 62 35 62 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 51 62 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 50 62 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 50 62 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 62 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 62 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 36 62 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 36 62 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 35 62 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 35 62 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 51 61 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 50 61 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 50 61 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 36 61 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 36 61 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 35 61 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 35 61 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 51 61 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 50 61 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 50 61 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 38 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 37 61 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 36 61 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 36 61 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 35 61 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 61 35 61 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 51 60 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 50 60 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 50 60 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 36 60 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 36 60 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 35 60 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 35 60 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 51 60 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 50 60 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 50 60 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 36 60 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 36 60 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 35 60 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 60 35 60 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 51 60 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 50 60 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 50 60 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 60 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 60 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 36 60 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 36 60 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 35 60 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 35 60 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 51 59 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 50 59 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 50 59 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 36 59 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 36 59 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 35 59 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 35 59 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 51 59 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 50 59 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 50 59 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 38 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 37 59 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 36 59 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 36 59 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 35 59 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 59 35 59 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 51 58 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 50 58 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 50 58 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 36 58 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 36 58 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 35 58 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 35 58 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 51 58 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 50 58 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 50 58 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 36 58 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 36 58 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 35 58 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 58 35 58 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 51 58 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 50 58 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 50 58 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 58 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 58 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 36 58 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 36 58 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 35 58 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 35 58 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 51 57 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 50 57 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 50 57 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 36 57 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 36 57 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 35 57 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 35 57 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 51 57 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 50 57 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 50 57 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 38 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 37 57 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 36 57 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 36 57 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 35 57 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 57 35 57 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 51 56 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 50 56 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 50 56 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 36 56 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 36 56 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 35 56 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 35 56 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 51 56 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 50 56 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 50 56 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 36 56 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 36 56 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 35 56 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 56 35 56 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 51 56 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 50 56 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 50 56 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 56 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 56 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 36 56 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 36 56 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 35 56 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 35 56 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 51 55 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 50 55 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 50 55 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 36 55 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 36 55 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 35 55 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 35 55 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 51 55 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 50 55 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 50 55 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 38 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 37 55 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 36 55 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 36 55 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 35 55 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 55 35 55 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 51 54 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 50 54 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 50 54 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 36 54 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 36 54 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 35 54 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 35 54 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 51 54 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 50 54 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 50 54 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 36 54 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 36 54 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 35 54 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 54 35 54 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 51 54 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 50 54 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 50 54 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 54 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 54 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 36 54 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 36 54 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 35 54 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 35 54 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 51 53 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 50 53 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 50 53 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 38 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 36 53 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 36 53 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 35 53 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 53 35 53 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 51 53 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 50 53 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 50 53 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 38 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 53 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 53 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 36 53 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 36 53 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 35 53 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 35 53 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 51 52 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 50 52 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 50 52 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 36 52 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 36 52 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 35 52 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 35 52 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 51 52 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 50 52 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 50 52 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 38 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 37 52 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 36 52 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 36 52 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 35 52 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 52 35 52 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 51 51 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 50 51 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 50 51 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 38 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 36 51 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 36 51 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 35 51 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 35 51 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 51 51 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 50 51 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 50 51 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 38 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 37 51 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 36 51 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 36 51 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 35 51 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 51 35 51 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 51 24 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 50 24 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 50 24 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 36 24 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 36 24 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 35 24 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 35 24 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 51 24 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 50 24 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 50 24 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 36 24 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 36 24 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 35 24 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 24 35 24 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 51 24 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 50 24 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 50 24 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 24 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 24 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 36 24 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 36 24 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 35 24 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 35 24 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 51 23 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 50 23 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 50 23 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 38 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 36 23 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 36 23 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 35 23 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 23 35 23 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 51 23 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 50 23 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 50 23 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 38 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 23 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 23 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 36 23 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 36 23 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 35 23 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 35 23 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 51 22 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 50 22 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 50 22 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 36 22 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 36 22 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 35 22 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 35 22 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 51 22 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 50 22 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 50 22 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 38 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 37 22 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 36 22 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 36 22 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 35 22 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 22 35 22 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 51 21 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 50 21 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 50 21 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 36 21 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 36 21 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 35 21 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 35 21 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 51 21 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 50 21 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 50 21 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 38 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 36 21 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 36 21 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 35 21 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 21 35 21 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 51 21 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 50 21 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 50 21 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 38 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 21 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 21 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 36 21 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 36 21 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 35 21 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 35 21 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 51 20 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 50 20 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 50 20 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 38 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 36 20 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 36 20 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 35 20 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 35 20 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 51 20 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 50 20 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 50 20 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 38 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 37 20 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 36 20 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 36 20 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 35 20 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 20 35 20 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 51 19 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 50 19 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 50 19 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 36 19 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 36 19 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 35 19 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 35 19 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 51 19 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 50 19 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 50 19 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 36 19 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 36 19 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 35 19 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 19 35 19 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 51 19 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 50 19 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 50 19 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 19 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 19 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 36 19 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 36 19 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 35 19 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 35 19 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 51 18 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 50 18 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 50 18 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 36 18 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 36 18 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 35 18 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 35 18 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 51 18 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 50 18 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 50 18 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 38 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 37 18 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 36 18 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 36 18 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 35 18 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 18 35 18 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 51 17 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 50 17 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 50 17 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 36 17 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 36 17 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 35 17 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 35 17 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 51 17 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 50 17 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 50 17 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 36 17 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 36 17 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 35 17 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 17 35 17 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 51 17 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 50 17 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 50 17 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 17 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 17 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 36 17 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 36 17 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 35 17 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 35 17 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 51 16 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 50 16 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 50 16 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 36 16 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 36 16 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 35 16 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 35 16 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 51 16 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 50 16 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 50 16 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 38 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 37 16 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 36 16 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 36 16 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 35 16 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 16 35 16 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 51 15 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 50 15 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 50 15 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 36 15 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 36 15 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 35 15 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 35 15 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 51 15 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 50 15 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 50 15 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 36 15 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 36 15 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 35 15 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 15 35 15 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 51 15 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 50 15 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 50 15 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 15 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 15 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 36 15 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 36 15 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 35 15 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 35 15 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 51 14 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 50 14 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 50 14 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 36 14 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 36 14 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 35 14 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 35 14 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 51 14 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 50 14 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 50 14 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 38 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 37 14 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 36 14 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 36 14 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 35 14 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 14 35 14 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 51 13 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 50 13 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 50 13 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 36 13 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 36 13 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 35 13 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 35 13 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 51 13 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 50 13 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 50 13 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 36 13 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 36 13 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 35 13 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 13 35 13 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 51 13 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 50 13 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 50 13 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 13 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 13 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 36 13 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 36 13 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 35 13 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 35 13 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 51 12 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 50 12 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 50 12 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 36 12 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 36 12 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 35 12 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 35 12 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 51 12 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 50 12 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 50 12 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 38 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 37 12 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 36 12 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 36 12 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 35 12 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 12 35 12 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 51 11 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 50 11 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 50 11 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 36 11 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 36 11 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 35 11 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 35 11 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 51 11 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 50 11 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 50 11 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 36 11 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 36 11 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 35 11 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 11 35 11 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 51 11 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 50 11 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 50 11 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 11 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 11 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 36 11 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 36 11 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 35 11 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 35 11 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 51 10 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 50 10 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 50 10 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 36 10 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 36 10 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 35 10 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 35 10 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 51 10 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 50 10 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 50 10 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 38 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 37 10 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 36 10 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 36 10 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 35 10 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 10 35 10 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 51 9 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 50 9 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 50 9 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 36 9 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 36 9 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 35 9 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 35 9 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 51 9 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 50 9 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 50 9 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 36 9 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 36 9 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 35 9 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 9 35 9 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 51 9 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 50 9 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 50 9 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 9 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 9 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 36 9 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 36 9 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 35 9 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 35 9 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 51 8 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 50 8 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 50 8 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 36 8 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 36 8 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 35 8 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 35 8 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 51 8 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 50 8 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 50 8 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 38 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 37 8 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 36 8 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 36 8 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 35 8 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 8 35 8 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 51 7 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 50 7 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 50 7 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 36 7 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 36 7 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 35 7 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 35 7 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 51 7 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 50 7 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 50 7 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 38 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 37 7 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 36 7 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 36 7 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 35 7 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 7 35 7 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 51 6 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 50 6 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 50 6 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 36 6 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 36 6 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 35 6 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 35 6 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 51 6 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 50 6 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 50 6 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 38 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 36 6 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 36 6 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 35 6 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 6 35 6 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 51 6 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 50 6 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 50 6 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 38 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 6 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 6 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 36 6 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 36 6 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 35 6 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 35 6 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 51 5 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 50 5 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 50 5 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 36 5 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 36 5 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 35 5 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 35 5 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 51 5 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 50 5 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 50 5 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 38 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 37 5 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 36 5 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 36 5 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 35 5 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 5 35 5 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 51 4 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 50 4 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 50 4 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 38 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 36 4 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 36 4 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 35 4 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 35 4 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 51 4 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 50 4 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 50 4 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 38 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 36 4 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 36 4 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 35 4 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 4 35 4 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 51 4 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 50 4 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 50 4 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 4 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 4 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 36 4 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 36 4 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 35 4 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 35 4 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 51 3 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 50 3 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 50 3 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 36 3 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 36 3 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 35 3 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 35 3 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 51 3 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 50 3 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 50 3 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 38 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 37 3 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 36 3 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 36 3 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 35 3 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 3 35 3 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 51 2 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 50 2 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 50 2 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 36 2 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 36 2 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 35 2 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 35 2 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 51 2 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 50 2 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 50 2 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 36 2 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 36 2 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 35 2 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 2 35 2 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 51 2 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 50 2 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 50 2 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 38 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 2 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 2 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 36 2 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 36 2 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 35 2 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 35 2 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 51 1 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 50 1 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 50 1 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 38 1 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 36 1 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 36 1 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 35 1 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 35 1 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 51 1 51 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 50 1 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 50 1 50 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 38 1 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 38 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 37 1 37 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 36 1 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 36 1 36 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 35 1 35 6 VSSA
port 8 nsew ground bidirectional
rlabel nfet_brown s 1 35 1 35 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 198
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
