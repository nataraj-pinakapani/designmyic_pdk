magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 2 3 3 6 DRAIN
port 1 nsew
rlabel rotate s 2 3 2 3 6 GATE
port 2 nsew
rlabel rotate s 2 3 2 3 6 GATE
port 2 nsew
rlabel rotate s 2 0 2 1 8 GATE
port 2 nsew
rlabel rotate s 2 0 2 0 8 GATE
port 2 nsew
rlabel rotate s 1 3 2 3 6 GATE
port 2 nsew
rlabel rotate s 1 3 2 3 6 GATE
port 2 nsew
rlabel rotate s 1 0 2 1 8 GATE
port 2 nsew
rlabel rotate s 1 0 2 0 8 GATE
port 2 nsew
rlabel  s 1 3 2 4 6 GATE
port 2 nsew
rlabel  s 1 0 2 1 8 GATE
port 2 nsew
rlabel  s 1 3 2 4 6 GATE
port 2 nsew
rlabel  s 1 0 2 1 8 GATE
port 2 nsew
rlabel  s 0 1 3 2 6 SOURCE
port 3 nsew
rlabel  s 0 1 1 3 4 SUBSTRATE
port 4 nsew
rlabel  s 3 1 3 3 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 3 4
string LEFview TRUE
<< end >>
