magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 0 0 976 1214
<< pmoslvt >>
rect 204 102 304 1112
rect 360 102 460 1112
rect 516 102 616 1112
rect 672 102 772 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 304 1100 360 1112
rect 304 1066 315 1100
rect 349 1066 360 1100
rect 304 1032 360 1066
rect 304 998 315 1032
rect 349 998 360 1032
rect 304 964 360 998
rect 304 930 315 964
rect 349 930 360 964
rect 304 896 360 930
rect 304 862 315 896
rect 349 862 360 896
rect 304 828 360 862
rect 304 794 315 828
rect 349 794 360 828
rect 304 760 360 794
rect 304 726 315 760
rect 349 726 360 760
rect 304 692 360 726
rect 304 658 315 692
rect 349 658 360 692
rect 304 624 360 658
rect 304 590 315 624
rect 349 590 360 624
rect 304 556 360 590
rect 304 522 315 556
rect 349 522 360 556
rect 304 488 360 522
rect 304 454 315 488
rect 349 454 360 488
rect 304 420 360 454
rect 304 386 315 420
rect 349 386 360 420
rect 304 352 360 386
rect 304 318 315 352
rect 349 318 360 352
rect 304 284 360 318
rect 304 250 315 284
rect 349 250 360 284
rect 304 216 360 250
rect 304 182 315 216
rect 349 182 360 216
rect 304 148 360 182
rect 304 114 315 148
rect 349 114 360 148
rect 304 102 360 114
rect 460 1100 516 1112
rect 460 1066 471 1100
rect 505 1066 516 1100
rect 460 1032 516 1066
rect 460 998 471 1032
rect 505 998 516 1032
rect 460 964 516 998
rect 460 930 471 964
rect 505 930 516 964
rect 460 896 516 930
rect 460 862 471 896
rect 505 862 516 896
rect 460 828 516 862
rect 460 794 471 828
rect 505 794 516 828
rect 460 760 516 794
rect 460 726 471 760
rect 505 726 516 760
rect 460 692 516 726
rect 460 658 471 692
rect 505 658 516 692
rect 460 624 516 658
rect 460 590 471 624
rect 505 590 516 624
rect 460 556 516 590
rect 460 522 471 556
rect 505 522 516 556
rect 460 488 516 522
rect 460 454 471 488
rect 505 454 516 488
rect 460 420 516 454
rect 460 386 471 420
rect 505 386 516 420
rect 460 352 516 386
rect 460 318 471 352
rect 505 318 516 352
rect 460 284 516 318
rect 460 250 471 284
rect 505 250 516 284
rect 460 216 516 250
rect 460 182 471 216
rect 505 182 516 216
rect 460 148 516 182
rect 460 114 471 148
rect 505 114 516 148
rect 460 102 516 114
rect 616 1100 672 1112
rect 616 1066 627 1100
rect 661 1066 672 1100
rect 616 1032 672 1066
rect 616 998 627 1032
rect 661 998 672 1032
rect 616 964 672 998
rect 616 930 627 964
rect 661 930 672 964
rect 616 896 672 930
rect 616 862 627 896
rect 661 862 672 896
rect 616 828 672 862
rect 616 794 627 828
rect 661 794 672 828
rect 616 760 672 794
rect 616 726 627 760
rect 661 726 672 760
rect 616 692 672 726
rect 616 658 627 692
rect 661 658 672 692
rect 616 624 672 658
rect 616 590 627 624
rect 661 590 672 624
rect 616 556 672 590
rect 616 522 627 556
rect 661 522 672 556
rect 616 488 672 522
rect 616 454 627 488
rect 661 454 672 488
rect 616 420 672 454
rect 616 386 627 420
rect 661 386 672 420
rect 616 352 672 386
rect 616 318 627 352
rect 661 318 672 352
rect 616 284 672 318
rect 616 250 627 284
rect 661 250 672 284
rect 616 216 672 250
rect 616 182 627 216
rect 661 182 672 216
rect 616 148 672 182
rect 616 114 627 148
rect 661 114 672 148
rect 616 102 672 114
rect 772 1100 828 1112
rect 772 1066 783 1100
rect 817 1066 828 1100
rect 772 1032 828 1066
rect 772 998 783 1032
rect 817 998 828 1032
rect 772 964 828 998
rect 772 930 783 964
rect 817 930 828 964
rect 772 896 828 930
rect 772 862 783 896
rect 817 862 828 896
rect 772 828 828 862
rect 772 794 783 828
rect 817 794 828 828
rect 772 760 828 794
rect 772 726 783 760
rect 817 726 828 760
rect 772 692 828 726
rect 772 658 783 692
rect 817 658 828 692
rect 772 624 828 658
rect 772 590 783 624
rect 817 590 828 624
rect 772 556 828 590
rect 772 522 783 556
rect 817 522 828 556
rect 772 488 828 522
rect 772 454 783 488
rect 817 454 828 488
rect 772 420 828 454
rect 772 386 783 420
rect 817 386 828 420
rect 772 352 828 386
rect 772 318 783 352
rect 817 318 828 352
rect 772 284 828 318
rect 772 250 783 284
rect 817 250 828 284
rect 772 216 828 250
rect 772 182 783 216
rect 817 182 828 216
rect 772 148 828 182
rect 772 114 783 148
rect 817 114 828 148
rect 772 102 828 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 315 1066 349 1100
rect 315 998 349 1032
rect 315 930 349 964
rect 315 862 349 896
rect 315 794 349 828
rect 315 726 349 760
rect 315 658 349 692
rect 315 590 349 624
rect 315 522 349 556
rect 315 454 349 488
rect 315 386 349 420
rect 315 318 349 352
rect 315 250 349 284
rect 315 182 349 216
rect 315 114 349 148
rect 471 1066 505 1100
rect 471 998 505 1032
rect 471 930 505 964
rect 471 862 505 896
rect 471 794 505 828
rect 471 726 505 760
rect 471 658 505 692
rect 471 590 505 624
rect 471 522 505 556
rect 471 454 505 488
rect 471 386 505 420
rect 471 318 505 352
rect 471 250 505 284
rect 471 182 505 216
rect 471 114 505 148
rect 627 1066 661 1100
rect 627 998 661 1032
rect 627 930 661 964
rect 627 862 661 896
rect 627 794 661 828
rect 627 726 661 760
rect 627 658 661 692
rect 627 590 661 624
rect 627 522 661 556
rect 627 454 661 488
rect 627 386 661 420
rect 627 318 661 352
rect 627 250 661 284
rect 627 182 661 216
rect 627 114 661 148
rect 783 1066 817 1100
rect 783 998 817 1032
rect 783 930 817 964
rect 783 862 817 896
rect 783 794 817 828
rect 783 726 817 760
rect 783 658 817 692
rect 783 590 817 624
rect 783 522 817 556
rect 783 454 817 488
rect 783 386 817 420
rect 783 318 817 352
rect 783 250 817 284
rect 783 182 817 216
rect 783 114 817 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 882 1066 940 1112
rect 882 1032 894 1066
rect 928 1032 940 1066
rect 882 998 940 1032
rect 882 964 894 998
rect 928 964 940 998
rect 882 930 940 964
rect 882 896 894 930
rect 928 896 940 930
rect 882 862 940 896
rect 882 828 894 862
rect 928 828 940 862
rect 882 794 940 828
rect 882 760 894 794
rect 928 760 940 794
rect 882 726 940 760
rect 882 692 894 726
rect 928 692 940 726
rect 882 658 940 692
rect 882 624 894 658
rect 928 624 940 658
rect 882 590 940 624
rect 882 556 894 590
rect 928 556 940 590
rect 882 522 940 556
rect 882 488 894 522
rect 928 488 940 522
rect 882 454 940 488
rect 882 420 894 454
rect 928 420 940 454
rect 882 386 940 420
rect 882 352 894 386
rect 928 352 940 386
rect 882 318 940 352
rect 882 284 894 318
rect 928 284 940 318
rect 882 250 940 284
rect 882 216 894 250
rect 928 216 940 250
rect 882 182 940 216
rect 882 148 894 182
rect 928 148 940 182
rect 882 102 940 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 894 1032 928 1066
rect 894 964 928 998
rect 894 896 928 930
rect 894 828 928 862
rect 894 760 928 794
rect 894 692 928 726
rect 894 624 928 658
rect 894 556 928 590
rect 894 488 928 522
rect 894 420 928 454
rect 894 352 928 386
rect 894 284 928 318
rect 894 216 928 250
rect 894 148 928 182
<< poly >>
rect 183 1194 793 1214
rect 183 1160 199 1194
rect 233 1160 267 1194
rect 301 1160 335 1194
rect 369 1160 403 1194
rect 437 1160 471 1194
rect 505 1160 539 1194
rect 573 1160 607 1194
rect 641 1160 675 1194
rect 709 1160 743 1194
rect 777 1160 793 1194
rect 183 1144 793 1160
rect 204 1112 304 1144
rect 360 1112 460 1144
rect 516 1112 616 1144
rect 672 1112 772 1144
rect 204 70 304 102
rect 360 70 460 102
rect 516 70 616 102
rect 672 70 772 102
rect 183 54 793 70
rect 183 20 199 54
rect 233 20 267 54
rect 301 20 335 54
rect 369 20 403 54
rect 437 20 471 54
rect 505 20 539 54
rect 573 20 607 54
rect 641 20 675 54
rect 709 20 743 54
rect 777 20 793 54
rect 183 0 793 20
<< polycont >>
rect 199 1160 233 1194
rect 267 1160 301 1194
rect 335 1160 369 1194
rect 403 1160 437 1194
rect 471 1160 505 1194
rect 539 1160 573 1194
rect 607 1160 641 1194
rect 675 1160 709 1194
rect 743 1160 777 1194
rect 199 20 233 54
rect 267 20 301 54
rect 335 20 369 54
rect 403 20 437 54
rect 471 20 505 54
rect 539 20 573 54
rect 607 20 641 54
rect 675 20 709 54
rect 743 20 777 54
<< locali >>
rect 233 1160 255 1194
rect 301 1160 327 1194
rect 369 1160 399 1194
rect 437 1160 471 1194
rect 505 1160 539 1194
rect 577 1160 607 1194
rect 649 1160 675 1194
rect 721 1160 743 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 315 1100 349 1116
rect 315 1032 349 1058
rect 315 964 349 986
rect 315 896 349 914
rect 315 828 349 842
rect 315 760 349 770
rect 315 692 349 698
rect 315 624 349 626
rect 315 588 349 590
rect 315 516 349 522
rect 315 444 349 454
rect 315 372 349 386
rect 315 300 349 318
rect 315 228 349 250
rect 315 156 349 182
rect 315 98 349 114
rect 471 1100 505 1116
rect 471 1032 505 1058
rect 471 964 505 986
rect 471 896 505 914
rect 471 828 505 842
rect 471 760 505 770
rect 471 692 505 698
rect 471 624 505 626
rect 471 588 505 590
rect 471 516 505 522
rect 471 444 505 454
rect 471 372 505 386
rect 471 300 505 318
rect 471 228 505 250
rect 471 156 505 182
rect 471 98 505 114
rect 627 1100 661 1116
rect 627 1032 661 1058
rect 627 964 661 986
rect 627 896 661 914
rect 627 828 661 842
rect 627 760 661 770
rect 627 692 661 698
rect 627 624 661 626
rect 627 588 661 590
rect 627 516 661 522
rect 627 444 661 454
rect 627 372 661 386
rect 627 300 661 318
rect 627 228 661 250
rect 627 156 661 182
rect 627 98 661 114
rect 783 1100 817 1116
rect 783 1032 817 1058
rect 783 964 817 986
rect 783 896 817 914
rect 783 828 817 842
rect 783 760 817 770
rect 783 692 817 698
rect 783 624 817 626
rect 783 588 817 590
rect 783 516 817 522
rect 783 444 817 454
rect 783 372 817 386
rect 783 300 817 318
rect 783 228 817 250
rect 783 156 817 182
rect 894 1020 928 1032
rect 894 948 928 964
rect 894 876 928 896
rect 894 804 928 828
rect 894 732 928 760
rect 894 660 928 692
rect 894 590 928 624
rect 894 522 928 554
rect 894 454 928 482
rect 894 386 928 410
rect 894 318 928 338
rect 894 250 928 266
rect 894 182 928 194
rect 783 98 817 114
rect 233 20 255 54
rect 301 20 327 54
rect 369 20 399 54
rect 437 20 471 54
rect 505 20 539 54
rect 577 20 607 54
rect 649 20 675 54
rect 721 20 743 54
<< viali >>
rect 183 1160 199 1194
rect 199 1160 217 1194
rect 255 1160 267 1194
rect 267 1160 289 1194
rect 327 1160 335 1194
rect 335 1160 361 1194
rect 399 1160 403 1194
rect 403 1160 433 1194
rect 471 1160 505 1194
rect 543 1160 573 1194
rect 573 1160 577 1194
rect 615 1160 641 1194
rect 641 1160 649 1194
rect 687 1160 709 1194
rect 709 1160 721 1194
rect 759 1160 777 1194
rect 777 1160 793 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 315 1066 349 1092
rect 315 1058 349 1066
rect 315 998 349 1020
rect 315 986 349 998
rect 315 930 349 948
rect 315 914 349 930
rect 315 862 349 876
rect 315 842 349 862
rect 315 794 349 804
rect 315 770 349 794
rect 315 726 349 732
rect 315 698 349 726
rect 315 658 349 660
rect 315 626 349 658
rect 315 556 349 588
rect 315 554 349 556
rect 315 488 349 516
rect 315 482 349 488
rect 315 420 349 444
rect 315 410 349 420
rect 315 352 349 372
rect 315 338 349 352
rect 315 284 349 300
rect 315 266 349 284
rect 315 216 349 228
rect 315 194 349 216
rect 315 148 349 156
rect 315 122 349 148
rect 471 1066 505 1092
rect 471 1058 505 1066
rect 471 998 505 1020
rect 471 986 505 998
rect 471 930 505 948
rect 471 914 505 930
rect 471 862 505 876
rect 471 842 505 862
rect 471 794 505 804
rect 471 770 505 794
rect 471 726 505 732
rect 471 698 505 726
rect 471 658 505 660
rect 471 626 505 658
rect 471 556 505 588
rect 471 554 505 556
rect 471 488 505 516
rect 471 482 505 488
rect 471 420 505 444
rect 471 410 505 420
rect 471 352 505 372
rect 471 338 505 352
rect 471 284 505 300
rect 471 266 505 284
rect 471 216 505 228
rect 471 194 505 216
rect 471 148 505 156
rect 471 122 505 148
rect 627 1066 661 1092
rect 627 1058 661 1066
rect 627 998 661 1020
rect 627 986 661 998
rect 627 930 661 948
rect 627 914 661 930
rect 627 862 661 876
rect 627 842 661 862
rect 627 794 661 804
rect 627 770 661 794
rect 627 726 661 732
rect 627 698 661 726
rect 627 658 661 660
rect 627 626 661 658
rect 627 556 661 588
rect 627 554 661 556
rect 627 488 661 516
rect 627 482 661 488
rect 627 420 661 444
rect 627 410 661 420
rect 627 352 661 372
rect 627 338 661 352
rect 627 284 661 300
rect 627 266 661 284
rect 627 216 661 228
rect 627 194 661 216
rect 627 148 661 156
rect 627 122 661 148
rect 783 1066 817 1092
rect 783 1058 817 1066
rect 783 998 817 1020
rect 783 986 817 998
rect 783 930 817 948
rect 783 914 817 930
rect 783 862 817 876
rect 783 842 817 862
rect 783 794 817 804
rect 783 770 817 794
rect 783 726 817 732
rect 783 698 817 726
rect 783 658 817 660
rect 783 626 817 658
rect 783 556 817 588
rect 783 554 817 556
rect 783 488 817 516
rect 783 482 817 488
rect 783 420 817 444
rect 783 410 817 420
rect 783 352 817 372
rect 783 338 817 352
rect 783 284 817 300
rect 783 266 817 284
rect 783 216 817 228
rect 783 194 817 216
rect 783 148 817 156
rect 783 122 817 148
rect 894 1066 928 1092
rect 894 1058 928 1066
rect 894 998 928 1020
rect 894 986 928 998
rect 894 930 928 948
rect 894 914 928 930
rect 894 862 928 876
rect 894 842 928 862
rect 894 794 928 804
rect 894 770 928 794
rect 894 726 928 732
rect 894 698 928 726
rect 894 658 928 660
rect 894 626 928 658
rect 894 556 928 588
rect 894 554 928 556
rect 894 488 928 516
rect 894 482 928 488
rect 894 420 928 444
rect 894 410 928 420
rect 894 352 928 372
rect 894 338 928 352
rect 894 284 928 300
rect 894 266 928 284
rect 894 216 928 228
rect 894 194 928 216
rect 894 148 928 156
rect 894 122 928 148
rect 183 20 199 54
rect 199 20 217 54
rect 255 20 267 54
rect 267 20 289 54
rect 327 20 335 54
rect 335 20 361 54
rect 399 20 403 54
rect 403 20 433 54
rect 471 20 505 54
rect 543 20 573 54
rect 573 20 577 54
rect 615 20 641 54
rect 641 20 649 54
rect 687 20 709 54
rect 709 20 721 54
rect 759 20 777 54
rect 777 20 793 54
<< metal1 >>
rect 171 1194 805 1214
rect 171 1160 183 1194
rect 217 1160 255 1194
rect 289 1160 327 1194
rect 361 1160 399 1194
rect 433 1160 471 1194
rect 505 1160 543 1194
rect 577 1160 615 1194
rect 649 1160 687 1194
rect 721 1160 759 1194
rect 793 1160 805 1194
rect 171 1148 805 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 306 1098 358 1104
rect 306 1034 358 1046
rect 306 970 358 982
rect 306 914 315 918
rect 349 914 358 918
rect 306 906 358 914
rect 306 842 315 854
rect 349 842 358 854
rect 306 778 315 790
rect 349 778 358 790
rect 306 714 315 726
rect 349 714 358 726
rect 306 660 358 662
rect 306 626 315 660
rect 349 626 358 660
rect 306 588 358 626
rect 306 554 315 588
rect 349 554 358 588
rect 306 516 358 554
rect 306 482 315 516
rect 349 482 358 516
rect 306 444 358 482
rect 306 410 315 444
rect 349 410 358 444
rect 306 372 358 410
rect 306 338 315 372
rect 349 338 358 372
rect 306 300 358 338
rect 306 266 315 300
rect 349 266 358 300
rect 306 228 358 266
rect 306 194 315 228
rect 349 194 358 228
rect 306 156 358 194
rect 306 122 315 156
rect 349 122 358 156
rect 306 110 358 122
rect 462 1092 514 1104
rect 462 1058 471 1092
rect 505 1058 514 1092
rect 462 1020 514 1058
rect 462 986 471 1020
rect 505 986 514 1020
rect 462 948 514 986
rect 462 914 471 948
rect 505 914 514 948
rect 462 876 514 914
rect 462 842 471 876
rect 505 842 514 876
rect 462 804 514 842
rect 462 770 471 804
rect 505 770 514 804
rect 462 732 514 770
rect 462 698 471 732
rect 505 698 514 732
rect 462 660 514 698
rect 462 626 471 660
rect 505 626 514 660
rect 462 588 514 626
rect 462 554 471 588
rect 505 554 514 588
rect 462 552 514 554
rect 462 488 471 500
rect 505 488 514 500
rect 462 424 471 436
rect 505 424 514 436
rect 462 360 471 372
rect 505 360 514 372
rect 462 300 514 308
rect 462 296 471 300
rect 505 296 514 300
rect 462 232 514 244
rect 462 168 514 180
rect 462 110 514 116
rect 618 1098 670 1104
rect 618 1034 670 1046
rect 618 970 670 982
rect 618 914 627 918
rect 661 914 670 918
rect 618 906 670 914
rect 618 842 627 854
rect 661 842 670 854
rect 618 778 627 790
rect 661 778 670 790
rect 618 714 627 726
rect 661 714 670 726
rect 618 660 670 662
rect 618 626 627 660
rect 661 626 670 660
rect 618 588 670 626
rect 618 554 627 588
rect 661 554 670 588
rect 618 516 670 554
rect 618 482 627 516
rect 661 482 670 516
rect 618 444 670 482
rect 618 410 627 444
rect 661 410 670 444
rect 618 372 670 410
rect 618 338 627 372
rect 661 338 670 372
rect 618 300 670 338
rect 618 266 627 300
rect 661 266 670 300
rect 618 228 670 266
rect 618 194 627 228
rect 661 194 670 228
rect 618 156 670 194
rect 618 122 627 156
rect 661 122 670 156
rect 618 110 670 122
rect 774 1092 826 1104
rect 774 1058 783 1092
rect 817 1058 826 1092
rect 774 1020 826 1058
rect 774 986 783 1020
rect 817 986 826 1020
rect 774 948 826 986
rect 774 914 783 948
rect 817 914 826 948
rect 774 876 826 914
rect 774 842 783 876
rect 817 842 826 876
rect 774 804 826 842
rect 774 770 783 804
rect 817 770 826 804
rect 774 732 826 770
rect 774 698 783 732
rect 817 698 826 732
rect 774 660 826 698
rect 774 626 783 660
rect 817 626 826 660
rect 774 588 826 626
rect 774 554 783 588
rect 817 554 826 588
rect 774 552 826 554
rect 774 488 783 500
rect 817 488 826 500
rect 774 424 783 436
rect 817 424 826 436
rect 774 360 783 372
rect 817 360 826 372
rect 774 300 826 308
rect 774 296 783 300
rect 817 296 826 300
rect 774 232 826 244
rect 774 168 826 180
rect 774 110 826 116
rect 882 1092 940 1104
rect 882 1058 894 1092
rect 928 1058 940 1092
rect 882 1020 940 1058
rect 882 986 894 1020
rect 928 986 940 1020
rect 882 948 940 986
rect 882 914 894 948
rect 928 914 940 948
rect 882 876 940 914
rect 882 842 894 876
rect 928 842 940 876
rect 882 804 940 842
rect 882 770 894 804
rect 928 770 940 804
rect 882 732 940 770
rect 882 698 894 732
rect 928 698 940 732
rect 882 660 940 698
rect 882 626 894 660
rect 928 626 940 660
rect 882 588 940 626
rect 882 554 894 588
rect 928 554 940 588
rect 882 516 940 554
rect 882 482 894 516
rect 928 482 940 516
rect 882 444 940 482
rect 882 410 894 444
rect 928 410 940 444
rect 882 372 940 410
rect 882 338 894 372
rect 928 338 940 372
rect 882 300 940 338
rect 882 266 894 300
rect 928 266 940 300
rect 882 228 940 266
rect 882 194 894 228
rect 928 194 940 228
rect 882 156 940 194
rect 882 122 894 156
rect 928 122 940 156
rect 882 110 940 122
rect 171 54 805 66
rect 171 20 183 54
rect 217 20 255 54
rect 289 20 327 54
rect 361 20 399 54
rect 433 20 471 54
rect 505 20 543 54
rect 577 20 615 54
rect 649 20 687 54
rect 721 20 759 54
rect 793 20 805 54
rect 171 0 805 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 306 1092 358 1098
rect 306 1058 315 1092
rect 315 1058 349 1092
rect 349 1058 358 1092
rect 306 1046 358 1058
rect 306 1020 358 1034
rect 306 986 315 1020
rect 315 986 349 1020
rect 349 986 358 1020
rect 306 982 358 986
rect 306 948 358 970
rect 306 918 315 948
rect 315 918 349 948
rect 349 918 358 948
rect 306 876 358 906
rect 306 854 315 876
rect 315 854 349 876
rect 349 854 358 876
rect 306 804 358 842
rect 306 790 315 804
rect 315 790 349 804
rect 349 790 358 804
rect 306 770 315 778
rect 315 770 349 778
rect 349 770 358 778
rect 306 732 358 770
rect 306 726 315 732
rect 315 726 349 732
rect 349 726 358 732
rect 306 698 315 714
rect 315 698 349 714
rect 349 698 358 714
rect 306 662 358 698
rect 462 516 514 552
rect 462 500 471 516
rect 471 500 505 516
rect 505 500 514 516
rect 462 482 471 488
rect 471 482 505 488
rect 505 482 514 488
rect 462 444 514 482
rect 462 436 471 444
rect 471 436 505 444
rect 505 436 514 444
rect 462 410 471 424
rect 471 410 505 424
rect 505 410 514 424
rect 462 372 514 410
rect 462 338 471 360
rect 471 338 505 360
rect 505 338 514 360
rect 462 308 514 338
rect 462 266 471 296
rect 471 266 505 296
rect 505 266 514 296
rect 462 244 514 266
rect 462 228 514 232
rect 462 194 471 228
rect 471 194 505 228
rect 505 194 514 228
rect 462 180 514 194
rect 462 156 514 168
rect 462 122 471 156
rect 471 122 505 156
rect 505 122 514 156
rect 462 116 514 122
rect 618 1092 670 1098
rect 618 1058 627 1092
rect 627 1058 661 1092
rect 661 1058 670 1092
rect 618 1046 670 1058
rect 618 1020 670 1034
rect 618 986 627 1020
rect 627 986 661 1020
rect 661 986 670 1020
rect 618 982 670 986
rect 618 948 670 970
rect 618 918 627 948
rect 627 918 661 948
rect 661 918 670 948
rect 618 876 670 906
rect 618 854 627 876
rect 627 854 661 876
rect 661 854 670 876
rect 618 804 670 842
rect 618 790 627 804
rect 627 790 661 804
rect 661 790 670 804
rect 618 770 627 778
rect 627 770 661 778
rect 661 770 670 778
rect 618 732 670 770
rect 618 726 627 732
rect 627 726 661 732
rect 661 726 670 732
rect 618 698 627 714
rect 627 698 661 714
rect 661 698 670 714
rect 618 662 670 698
rect 774 516 826 552
rect 774 500 783 516
rect 783 500 817 516
rect 817 500 826 516
rect 774 482 783 488
rect 783 482 817 488
rect 817 482 826 488
rect 774 444 826 482
rect 774 436 783 444
rect 783 436 817 444
rect 817 436 826 444
rect 774 410 783 424
rect 783 410 817 424
rect 817 410 826 424
rect 774 372 826 410
rect 774 338 783 360
rect 783 338 817 360
rect 817 338 826 360
rect 774 308 826 338
rect 774 266 783 296
rect 783 266 817 296
rect 817 266 826 296
rect 774 244 826 266
rect 774 228 826 232
rect 774 194 783 228
rect 783 194 817 228
rect 817 194 826 228
rect 774 180 826 194
rect 774 156 826 168
rect 774 122 783 156
rect 783 122 817 156
rect 817 122 826 156
rect 774 116 826 122
<< metal2 >>
rect 10 1098 966 1104
rect 10 1046 306 1098
rect 358 1046 618 1098
rect 670 1046 966 1098
rect 10 1034 966 1046
rect 10 982 306 1034
rect 358 982 618 1034
rect 670 982 966 1034
rect 10 970 966 982
rect 10 918 306 970
rect 358 918 618 970
rect 670 918 966 970
rect 10 906 966 918
rect 10 854 306 906
rect 358 854 618 906
rect 670 854 966 906
rect 10 842 966 854
rect 10 790 306 842
rect 358 790 618 842
rect 670 790 966 842
rect 10 778 966 790
rect 10 726 306 778
rect 358 726 618 778
rect 670 726 966 778
rect 10 714 966 726
rect 10 662 306 714
rect 358 662 618 714
rect 670 662 966 714
rect 10 632 966 662
rect 10 552 966 582
rect 10 500 150 552
rect 202 500 462 552
rect 514 500 774 552
rect 826 500 966 552
rect 10 488 966 500
rect 10 436 150 488
rect 202 436 462 488
rect 514 436 774 488
rect 826 436 966 488
rect 10 424 966 436
rect 10 372 150 424
rect 202 372 462 424
rect 514 372 774 424
rect 826 372 966 424
rect 10 360 966 372
rect 10 308 150 360
rect 202 308 462 360
rect 514 308 774 360
rect 826 308 966 360
rect 10 296 966 308
rect 10 244 150 296
rect 202 244 462 296
rect 514 244 774 296
rect 826 244 966 296
rect 10 232 966 244
rect 10 180 150 232
rect 202 180 462 232
rect 514 180 774 232
rect 826 180 966 232
rect 10 168 966 180
rect 10 116 150 168
rect 202 116 462 168
rect 514 116 774 168
rect 826 116 966 168
rect 10 110 966 116
<< labels >>
flabel metal2 s 13 771 32 841 0 FreeSans 400 90 0 0 DRAIN
port 1 nsew
flabel metal2 s 16 300 37 364 0 FreeSans 400 90 0 0 SOURCE
port 2 nsew
flabel metal1 s 58 732 58 732 7 FreeSans 400 90 0 0 BULK
port 3 nsew
flabel metal1 s 908 732 908 732 7 FreeSans 400 90 0 0 BULK
port 3 nsew
flabel metal1 s 171 1148 805 1214 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 171 0 805 66 0 FreeSans 300 0 0 0 GATE
port 4 nsew
<< properties >>
string GDS_END 10051678
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 10029198
<< end >>
