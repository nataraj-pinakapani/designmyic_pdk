/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/sky130_fd_pr__cap_var_hvt_fail.cdl