magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 53 75 56 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 48 75 51 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 9 1 14 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 9 75 14 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 9 1 13 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 9 75 13 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 69 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 64 1 68 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 68 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 1 48 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 52 1 53 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 56 1 57 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 48 75 48 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 52 75 53 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 56 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 1 57 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 48 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 1 42 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel 
 s 50 42 74 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 42 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 50 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 46 74 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 46 74 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 45 74 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 45 74 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 46 74 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 46 74 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 45 74 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 45 74 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 46 73 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 46 73 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 45 73 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 45 73 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 46 73 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 46 73 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 45 73 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 45 73 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 46 73 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 46 73 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 45 73 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 45 73 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 46 72 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 46 72 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 45 72 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 45 72 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 46 72 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 46 72 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 45 72 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 45 72 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 46 71 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 46 71 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 45 71 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 45 71 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 46 71 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 46 71 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 45 71 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 45 71 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 46 71 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 46 71 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 45 71 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 45 71 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 46 70 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 46 70 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 45 70 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 45 70 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 46 70 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 46 70 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 45 70 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 45 70 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 46 69 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 46 69 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 45 69 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 45 69 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 46 69 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 46 69 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 45 69 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 45 69 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 46 69 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 46 69 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 45 69 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 45 69 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 46 68 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 46 68 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 45 68 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 45 68 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 46 68 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 46 68 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 45 68 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 45 68 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 46 67 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 46 67 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 45 67 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 45 67 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 46 67 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 46 67 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 45 67 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 45 67 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 46 67 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 46 67 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 45 67 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 45 67 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 46 66 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 46 66 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 45 66 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 45 66 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 46 66 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 46 66 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 45 66 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 45 66 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 46 65 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 46 65 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 45 65 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 45 65 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 46 65 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 46 65 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 45 65 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 45 65 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 46 64 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 46 64 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 45 64 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 45 64 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 46 64 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 46 64 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 45 64 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 45 64 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 46 64 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 46 64 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 45 64 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 45 64 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 46 63 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 46 63 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 45 63 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 45 63 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 46 63 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 46 63 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 45 63 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 45 63 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 46 62 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 46 62 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 45 62 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 45 62 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 46 62 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 46 62 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 45 62 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 45 62 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 46 62 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 46 62 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 45 62 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 45 62 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 46 61 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 46 61 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 45 61 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 45 61 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 46 61 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 46 61 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 45 61 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 45 61 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 46 60 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 46 60 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 45 60 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 45 60 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 46 60 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 46 60 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 45 60 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 45 60 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 46 60 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 46 60 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 45 60 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 45 60 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 46 59 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 46 59 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 45 59 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 45 59 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 46 59 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 46 59 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 45 59 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 45 59 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 46 58 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 46 58 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 45 58 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 45 58 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 46 58 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 46 58 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 45 58 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 45 58 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 46 58 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 46 58 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 45 58 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 45 58 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 46 57 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 46 57 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 45 57 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 45 57 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 46 57 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 46 57 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 45 57 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 45 57 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 46 56 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 46 56 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 45 56 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 45 56 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 46 56 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 46 56 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 45 56 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 45 56 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 46 56 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 46 56 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 45 56 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 45 56 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 46 55 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 46 55 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 45 55 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 45 55 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 46 55 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 46 55 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 45 55 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 45 55 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 46 54 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 46 54 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 45 54 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 45 54 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 46 54 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 46 54 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 45 54 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 45 54 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 46 54 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 46 54 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 45 54 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 45 54 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 46 53 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 46 53 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 45 53 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 45 53 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 46 53 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 46 53 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 45 53 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 45 53 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 46 52 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 46 52 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 45 52 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 45 52 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 46 52 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 46 52 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 45 52 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 45 52 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 46 52 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 46 52 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 45 52 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 45 52 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 46 51 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 46 51 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 45 51 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 45 51 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 46 51 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 46 51 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 45 51 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 45 51 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 43 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 50 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 46 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 46 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 45 24 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 45 24 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 46 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 46 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 45 24 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 45 24 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 46 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 46 24 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 45 24 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 45 24 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 46 23 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 46 23 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 45 23 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 45 23 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 46 23 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 46 23 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 45 23 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 45 23 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 46 22 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 46 22 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 45 22 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 45 22 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 46 22 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 46 22 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 45 22 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 45 22 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 46 22 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 46 22 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 45 22 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 45 22 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 46 21 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 46 21 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 45 21 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 45 21 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 46 21 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 46 21 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 45 21 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 45 21 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 46 20 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 46 20 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 45 20 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 45 20 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 46 20 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 46 20 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 45 20 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 45 20 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 46 19 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 46 19 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 45 19 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 45 19 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 46 19 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 46 19 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 45 19 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 45 19 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 46 19 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 46 19 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 45 19 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 45 19 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 46 18 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 46 18 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 45 18 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 45 18 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 46 18 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 46 18 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 45 18 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 45 18 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 46 17 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 46 17 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 45 17 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 45 17 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 46 17 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 46 17 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 45 17 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 45 17 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 46 17 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 46 17 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 45 17 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 45 17 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 46 16 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 46 16 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 45 16 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 45 16 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 46 16 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 46 16 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 45 16 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 45 16 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 46 15 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 46 15 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 45 15 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 45 15 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 46 15 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 46 15 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 45 15 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 45 15 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 46 15 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 46 15 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 45 15 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 45 15 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 46 14 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 46 14 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 45 14 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 45 14 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 46 14 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 46 14 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 45 14 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 45 14 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 46 13 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 46 13 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 45 13 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 45 13 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 46 13 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 46 13 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 45 13 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 45 13 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 46 13 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 46 13 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 45 13 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 45 13 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 46 12 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 46 12 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 45 12 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 45 12 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 46 12 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 46 12 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 45 12 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 45 12 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 46 11 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 46 11 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 45 11 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 45 11 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 46 11 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 46 11 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 45 11 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 45 11 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 46 11 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 46 11 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 45 11 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 45 11 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 46 10 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 46 10 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 45 10 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 45 10 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 46 10 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 46 10 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 45 10 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 45 10 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 46 9 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 46 9 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 45 9 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 45 9 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 46 9 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 46 9 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 45 9 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 45 9 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 46 9 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 46 9 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 45 9 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 45 9 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 46 8 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 46 8 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 45 8 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 45 8 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 46 8 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 46 8 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 45 8 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 45 8 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 46 7 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 46 7 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 45 7 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 45 7 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 46 7 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 46 7 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 45 7 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 45 7 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 46 7 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 46 7 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 45 7 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 45 7 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 46 6 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 46 6 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 45 6 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 45 6 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 46 6 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 46 6 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 45 6 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 45 6 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 46 5 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 46 5 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 45 5 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 45 5 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 46 5 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 46 5 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 45 5 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 45 5 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 46 5 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 46 5 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 45 5 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 45 5 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 46 4 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 46 4 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 45 4 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 45 4 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 46 4 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 46 4 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 45 4 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 45 4 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 46 3 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 46 3 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 45 3 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 45 3 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 46 3 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 46 3 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 45 3 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 45 3 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 46 2 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 46 2 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 45 2 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 45 2 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 46 2 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 46 2 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 45 2 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 45 2 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 46 2 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 46 2 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 45 2 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 45 2 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 46 1 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 46 1 46 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 45 1 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 45 1 45 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 1 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 1 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 1 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 1 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 1 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
