magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 48 735 201
rect 0 0 736 48
<< scnmos >>
rect 79 47 109 175
rect 151 47 181 175
rect 363 47 393 175
rect 435 47 465 175
rect 531 47 561 175
rect 627 47 657 175
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 363 297 393 497
rect 447 297 477 497
rect 531 297 561 497
rect 627 297 657 497
<< ndiff >>
rect 27 161 79 175
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 47 151 175
rect 181 93 363 175
rect 181 59 191 93
rect 225 59 259 93
rect 293 59 363 93
rect 181 47 363 59
rect 393 47 435 175
rect 465 163 531 175
rect 465 129 479 163
rect 513 129 531 163
rect 465 93 531 129
rect 465 59 479 93
rect 513 59 531 93
rect 465 47 531 59
rect 561 47 627 175
rect 657 161 709 175
rect 657 127 667 161
rect 701 127 709 161
rect 657 93 709 127
rect 657 59 667 93
rect 701 59 709 93
rect 657 47 709 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 416 79 451
rect 27 382 35 416
rect 69 382 79 416
rect 27 347 79 382
rect 27 313 35 347
rect 69 313 79 347
rect 27 297 79 313
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 350 245 497
rect 193 316 203 350
rect 237 316 245 350
rect 193 297 245 316
rect 311 399 363 497
rect 311 365 319 399
rect 353 365 363 399
rect 311 297 363 365
rect 393 477 447 497
rect 393 443 403 477
rect 437 443 447 477
rect 393 297 447 443
rect 477 485 531 497
rect 477 451 487 485
rect 521 451 531 485
rect 477 416 531 451
rect 477 382 487 416
rect 521 382 531 416
rect 477 347 531 382
rect 477 313 487 347
rect 521 313 531 347
rect 477 297 531 313
rect 561 485 627 497
rect 561 451 571 485
rect 605 451 627 485
rect 561 415 627 451
rect 561 381 571 415
rect 605 381 627 415
rect 561 297 627 381
rect 657 485 709 497
rect 657 451 667 485
rect 701 451 709 485
rect 657 416 709 451
rect 657 382 667 416
rect 701 382 709 416
rect 657 347 709 382
rect 657 313 667 347
rect 701 313 709 347
rect 657 297 709 313
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 191 59 225 93
rect 259 59 293 93
rect 479 129 513 163
rect 479 59 513 93
rect 667 127 701 161
rect 667 59 701 93
<< pdiffc >>
rect 35 451 69 485
rect 35 382 69 416
rect 35 313 69 347
rect 119 443 153 477
rect 119 375 153 409
rect 203 316 237 350
rect 319 365 353 399
rect 403 443 437 477
rect 487 451 521 485
rect 487 382 521 416
rect 487 313 521 347
rect 571 451 605 485
rect 571 381 605 415
rect 667 451 701 485
rect 667 382 701 416
rect 667 313 701 347
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 363 497 393 523
rect 447 497 477 523
rect 531 497 561 523
rect 627 497 657 523
rect 79 266 109 297
rect 163 266 193 297
rect 363 266 393 297
rect 447 266 477 297
rect 531 266 561 297
rect 627 266 657 297
rect 21 250 109 266
rect 21 216 59 250
rect 93 216 109 250
rect 21 200 109 216
rect 79 175 109 200
rect 151 250 205 266
rect 151 216 161 250
rect 195 216 205 250
rect 151 200 205 216
rect 331 250 393 266
rect 331 216 347 250
rect 381 216 393 250
rect 331 200 393 216
rect 151 175 181 200
rect 363 175 393 200
rect 435 250 489 266
rect 435 216 445 250
rect 479 216 489 250
rect 435 200 489 216
rect 531 250 585 266
rect 531 216 541 250
rect 575 216 585 250
rect 531 200 585 216
rect 627 250 681 266
rect 627 216 637 250
rect 671 216 681 250
rect 627 200 681 216
rect 435 175 465 200
rect 531 175 561 200
rect 627 175 657 200
rect 79 21 109 47
rect 151 21 181 47
rect 363 21 393 47
rect 435 21 465 47
rect 531 21 561 47
rect 627 21 657 47
<< polycont >>
rect 59 216 93 250
rect 161 216 195 250
rect 347 216 381 250
rect 445 216 479 250
rect 541 216 575 250
rect 637 216 671 250
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 485 85 493
rect 19 451 35 485
rect 69 451 85 485
rect 119 477 437 493
rect 19 416 69 451
rect 19 382 35 416
rect 153 459 403 477
rect 119 415 153 443
rect 403 427 437 443
rect 471 485 537 493
rect 471 451 487 485
rect 521 451 537 485
rect 571 485 605 527
rect 651 485 719 493
rect 651 451 667 485
rect 701 451 719 485
rect 471 416 521 451
rect 19 347 69 382
rect 103 409 169 415
rect 103 375 119 409
rect 153 375 169 409
rect 19 313 35 347
rect 203 350 237 366
rect 303 365 319 399
rect 353 396 383 399
rect 353 394 387 396
rect 353 393 394 394
rect 353 365 403 393
rect 471 382 487 416
rect 571 415 605 451
rect 667 416 719 451
rect 471 365 521 382
rect 555 381 571 415
rect 605 381 621 415
rect 701 382 719 416
rect 69 334 85 336
rect 69 316 203 334
rect 369 347 521 365
rect 667 347 719 382
rect 237 316 285 334
rect 369 331 487 347
rect 69 313 285 316
rect 19 300 285 313
rect 471 313 487 331
rect 521 334 537 347
rect 644 334 667 347
rect 521 313 667 334
rect 701 313 719 347
rect 471 300 719 313
rect 19 297 85 300
rect 251 266 285 300
rect 17 250 109 263
rect 17 216 59 250
rect 93 216 109 250
rect 17 200 109 216
rect 143 250 217 263
rect 143 216 161 250
rect 195 216 217 250
rect 143 200 217 216
rect 251 163 296 266
rect 331 250 393 266
rect 331 216 347 250
rect 381 216 393 250
rect 331 200 393 216
rect 427 250 489 266
rect 427 216 445 250
rect 479 216 489 250
rect 427 200 489 216
rect 523 250 585 266
rect 523 216 541 250
rect 575 216 585 250
rect 523 200 585 216
rect 619 250 687 266
rect 619 216 637 250
rect 671 216 687 250
rect 619 200 687 216
rect 19 161 479 163
rect 19 127 35 161
rect 69 129 479 161
rect 513 129 529 163
rect 69 127 85 129
rect 19 93 85 127
rect 463 93 529 129
rect 19 59 35 93
rect 69 59 85 93
rect 19 51 85 59
rect 175 59 191 93
rect 225 59 259 93
rect 293 59 321 93
rect 463 59 479 93
rect 513 59 529 93
rect 651 161 717 163
rect 651 127 667 161
rect 701 127 717 161
rect 651 93 717 127
rect 651 59 667 93
rect 701 59 717 93
rect 175 17 321 59
rect 651 17 717 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a222oi_1
flabel pwell s 0 0 736 48 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 496 736 544 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
flabel metal1 s 0 496 736 544 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel metal1 s 0 0 736 48 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel locali s 164 218 198 252 0 FreeSans 340 0 0 0 C2
port 6 nsew signal input
flabel locali s 31 218 65 252 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 445 218 479 252 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 643 214 677 248 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 541 218 575 252 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 251 218 285 252 0 FreeSans 340 0 0 0 Y
port 11 nsew signal output
flabel locali s 351 218 385 252 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 736 48 1 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3694874
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3687786
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
