magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 831 47 861 177
rect 915 47 945 177
rect 1111 47 1141 177
rect 1195 47 1225 177
rect 1279 47 1309 177
rect 1363 47 1393 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 519 297 549 497
rect 603 297 633 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 939 297 969 497
rect 1035 297 1065 497
rect 1119 297 1149 497
rect 1279 297 1309 497
rect 1363 297 1393 497
<< ndiff >>
rect 27 97 79 177
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 93 163 127
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 161 331 177
rect 277 127 287 161
rect 321 127 331 161
rect 277 93 331 127
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 93 415 177
rect 361 59 371 93
rect 405 59 415 93
rect 361 47 415 59
rect 445 161 503 177
rect 445 127 459 161
rect 493 127 503 161
rect 445 93 503 127
rect 445 59 459 93
rect 493 59 503 93
rect 445 47 503 59
rect 533 93 587 177
rect 533 59 543 93
rect 577 59 587 93
rect 533 47 587 59
rect 617 161 671 177
rect 617 127 627 161
rect 661 127 671 161
rect 617 93 671 127
rect 617 59 627 93
rect 661 59 671 93
rect 617 47 671 59
rect 701 93 831 177
rect 701 59 711 93
rect 745 59 779 93
rect 813 59 831 93
rect 701 47 831 59
rect 861 161 915 177
rect 861 127 871 161
rect 905 127 915 161
rect 861 93 915 127
rect 861 59 871 93
rect 905 59 915 93
rect 861 47 915 59
rect 945 93 997 177
rect 945 59 955 93
rect 989 59 997 93
rect 945 47 997 59
rect 1059 93 1111 177
rect 1059 59 1067 93
rect 1101 59 1111 93
rect 1059 47 1111 59
rect 1141 163 1195 177
rect 1141 129 1151 163
rect 1185 129 1195 163
rect 1141 47 1195 129
rect 1225 161 1279 177
rect 1225 127 1235 161
rect 1269 127 1279 161
rect 1225 93 1279 127
rect 1225 59 1235 93
rect 1269 59 1279 93
rect 1225 47 1279 59
rect 1309 165 1363 177
rect 1309 131 1319 165
rect 1353 131 1363 165
rect 1309 47 1363 131
rect 1393 165 1445 177
rect 1393 131 1403 165
rect 1437 131 1445 165
rect 1393 93 1445 131
rect 1393 59 1403 93
rect 1437 59 1445 93
rect 1393 47 1445 59
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 425 163 497
rect 109 391 119 425
rect 153 391 163 425
rect 109 357 163 391
rect 109 323 119 357
rect 153 323 163 357
rect 109 297 163 323
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 409 331 497
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 477 413 497
rect 361 443 371 477
rect 405 443 413 477
rect 361 409 413 443
rect 361 375 371 409
rect 405 375 413 409
rect 361 297 413 375
rect 467 485 519 497
rect 467 451 475 485
rect 509 451 519 485
rect 467 297 519 451
rect 549 343 603 497
rect 549 309 559 343
rect 593 309 603 343
rect 549 297 603 309
rect 633 485 687 497
rect 633 451 643 485
rect 677 451 687 485
rect 633 297 687 451
rect 717 343 771 497
rect 717 309 727 343
rect 761 309 771 343
rect 717 297 771 309
rect 801 485 855 497
rect 801 451 811 485
rect 845 451 855 485
rect 801 297 855 451
rect 885 477 939 497
rect 885 443 895 477
rect 929 443 939 477
rect 885 409 939 443
rect 885 375 895 409
rect 929 375 939 409
rect 885 297 939 375
rect 969 485 1035 497
rect 969 451 979 485
rect 1013 451 1035 485
rect 969 297 1035 451
rect 1065 477 1119 497
rect 1065 443 1075 477
rect 1109 443 1119 477
rect 1065 409 1119 443
rect 1065 375 1075 409
rect 1109 375 1119 409
rect 1065 297 1119 375
rect 1149 485 1279 497
rect 1149 451 1159 485
rect 1193 451 1279 485
rect 1149 297 1279 451
rect 1309 477 1363 497
rect 1309 443 1319 477
rect 1353 443 1363 477
rect 1309 409 1363 443
rect 1309 375 1319 409
rect 1353 375 1363 409
rect 1309 297 1363 375
rect 1393 485 1445 497
rect 1393 451 1403 485
rect 1437 451 1445 485
rect 1393 393 1445 451
rect 1393 359 1403 393
rect 1437 359 1445 393
rect 1393 297 1445 359
<< ndiffc >>
rect 35 63 69 97
rect 119 127 153 161
rect 119 59 153 93
rect 203 59 237 93
rect 287 127 321 161
rect 287 59 321 93
rect 371 59 405 93
rect 459 127 493 161
rect 459 59 493 93
rect 543 59 577 93
rect 627 127 661 161
rect 627 59 661 93
rect 711 59 745 93
rect 779 59 813 93
rect 871 127 905 161
rect 871 59 905 93
rect 955 59 989 93
rect 1067 59 1101 93
rect 1151 129 1185 163
rect 1235 127 1269 161
rect 1235 59 1269 93
rect 1319 131 1353 165
rect 1403 131 1437 165
rect 1403 59 1437 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 391 153 425
rect 119 323 153 357
rect 203 443 237 477
rect 203 375 237 409
rect 287 375 321 409
rect 371 443 405 477
rect 371 375 405 409
rect 475 451 509 485
rect 559 309 593 343
rect 643 451 677 485
rect 727 309 761 343
rect 811 451 845 485
rect 895 443 929 477
rect 895 375 929 409
rect 979 451 1013 485
rect 1075 443 1109 477
rect 1075 375 1109 409
rect 1159 451 1193 485
rect 1319 443 1353 477
rect 1319 375 1353 409
rect 1403 451 1437 485
rect 1403 359 1437 393
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 519 497 549 523
rect 603 497 633 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 939 497 969 523
rect 1035 497 1065 523
rect 1119 497 1149 523
rect 1279 497 1309 523
rect 1363 497 1393 523
rect 79 265 109 297
rect 163 265 193 297
rect 22 249 193 265
rect 247 259 277 297
rect 331 259 361 297
rect 519 259 549 297
rect 603 259 633 297
rect 687 282 717 297
rect 771 282 801 297
rect 687 259 801 282
rect 22 215 32 249
rect 66 215 193 249
rect 22 199 193 215
rect 79 177 109 199
rect 163 177 193 199
rect 235 249 361 259
rect 235 215 251 249
rect 285 215 361 249
rect 235 195 361 215
rect 403 252 801 259
rect 855 282 885 297
rect 939 282 969 297
rect 403 249 789 252
rect 403 215 419 249
rect 453 215 491 249
rect 525 215 671 249
rect 705 215 739 249
rect 773 215 789 249
rect 855 249 969 282
rect 855 222 919 249
rect 403 205 789 215
rect 831 215 919 222
rect 953 215 969 249
rect 247 177 277 195
rect 331 177 361 195
rect 415 177 445 205
rect 503 199 701 205
rect 503 177 533 199
rect 587 177 617 199
rect 671 177 701 199
rect 831 192 969 215
rect 1035 259 1065 297
rect 1119 259 1149 297
rect 1279 265 1309 297
rect 1363 265 1393 297
rect 1035 249 1225 259
rect 1035 215 1067 249
rect 1101 215 1158 249
rect 1192 215 1225 249
rect 1035 205 1225 215
rect 831 177 861 192
rect 915 177 945 192
rect 1111 177 1141 205
rect 1195 177 1225 205
rect 1279 249 1451 265
rect 1279 215 1405 249
rect 1439 215 1451 249
rect 1279 199 1451 215
rect 1279 177 1309 199
rect 1363 177 1393 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
rect 831 21 861 47
rect 915 21 945 47
rect 1111 21 1141 47
rect 1195 21 1225 47
rect 1279 21 1309 47
rect 1363 21 1393 47
<< polycont >>
rect 32 215 66 249
rect 251 215 285 249
rect 419 215 453 249
rect 491 215 525 249
rect 671 215 705 249
rect 739 215 773 249
rect 919 215 953 249
rect 1067 215 1101 249
rect 1158 215 1192 249
rect 1405 215 1439 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 35 477 405 493
rect 69 459 203 477
rect 35 409 69 443
rect 237 459 371 477
rect 103 391 119 425
rect 153 391 169 425
rect 203 409 237 443
rect 459 485 525 527
rect 459 451 475 485
rect 509 451 525 485
rect 627 485 693 527
rect 627 451 643 485
rect 677 451 693 485
rect 795 485 861 527
rect 795 451 811 485
rect 845 451 861 485
rect 895 477 929 493
rect 35 359 69 375
rect 119 357 153 391
rect 203 359 237 375
rect 287 409 321 425
rect 27 249 70 325
rect 27 215 32 249
rect 66 215 70 249
rect 27 149 70 215
rect 287 325 321 375
rect 371 409 405 443
rect 963 485 1035 527
rect 963 451 979 485
rect 1013 451 1035 485
rect 1075 477 1109 493
rect 895 417 929 443
rect 1143 485 1209 527
rect 1143 451 1159 485
rect 1193 451 1209 485
rect 1319 477 1353 493
rect 1075 417 1109 443
rect 1319 417 1353 443
rect 371 359 405 375
rect 439 409 1353 417
rect 439 383 895 409
rect 439 325 477 383
rect 929 383 1075 409
rect 895 359 929 375
rect 1109 383 1319 409
rect 1075 359 1109 375
rect 1319 359 1353 375
rect 1387 485 1454 527
rect 1387 451 1403 485
rect 1437 451 1454 485
rect 1387 393 1454 451
rect 1387 359 1403 393
rect 1437 359 1454 393
rect 119 177 153 323
rect 212 257 251 325
rect 287 291 477 325
rect 543 309 559 343
rect 593 309 727 343
rect 761 309 777 343
rect 212 249 301 257
rect 212 215 251 249
rect 285 215 301 249
rect 371 215 419 249
rect 453 215 491 249
rect 525 215 541 249
rect 371 177 405 215
rect 582 177 621 309
rect 830 291 1337 325
rect 830 249 864 291
rect 655 215 671 249
rect 705 215 739 249
rect 773 215 864 249
rect 903 249 989 257
rect 903 215 919 249
rect 953 215 989 249
rect 1051 249 1208 257
rect 1051 215 1067 249
rect 1101 215 1158 249
rect 1192 215 1208 249
rect 119 161 405 177
rect 153 143 287 161
rect 19 97 69 113
rect 19 63 35 97
rect 119 93 153 127
rect 321 143 405 161
rect 459 161 661 177
rect 203 93 237 109
rect 287 93 321 127
rect 493 143 627 161
rect 371 93 405 109
rect 459 93 493 127
rect 543 93 577 109
rect 627 93 661 127
rect 871 163 1201 177
rect 871 161 1151 163
rect 905 143 1151 161
rect 1135 129 1151 143
rect 1185 129 1201 163
rect 1235 161 1269 177
rect 711 93 813 109
rect 871 93 905 127
rect 1303 165 1337 291
rect 1389 249 1455 323
rect 1389 215 1405 249
rect 1439 215 1455 249
rect 1403 165 1454 181
rect 1303 131 1319 165
rect 1353 131 1369 165
rect 1303 129 1369 131
rect 1437 131 1454 165
rect 955 93 989 109
rect 1235 93 1269 127
rect 1403 100 1454 131
rect 19 17 69 63
rect 103 59 119 93
rect 153 59 169 93
rect 271 59 287 93
rect 321 59 337 93
rect 439 59 459 93
rect 493 59 509 93
rect 611 59 627 93
rect 661 59 677 93
rect 745 59 779 93
rect 855 59 871 93
rect 905 59 921 93
rect 203 17 237 59
rect 371 17 405 59
rect 543 17 577 59
rect 711 17 813 59
rect 955 17 989 59
rect 1051 59 1067 93
rect 1101 59 1235 93
rect 1387 93 1454 100
rect 1387 85 1403 93
rect 1269 59 1403 85
rect 1437 59 1454 93
rect 1051 51 1454 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1409 221 1443 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 1150 221 1184 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1058 221 1092 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 586 153 620 187 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 586 289 620 323 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
rlabel comment s 0 0 0 0 4 a311o_4
flabel comment s 556 227 556 227 0 FreeSans 200 0 0 0 no_jumper_check
rlabel metal1 s 0 -48 1472 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 3720592
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3708870
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 36.800 0.000 
<< end >>
