magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 11 0 11 12 6 C0
port 1 nsew
rlabel  s 9 6 10 11 6 C0
port 1 nsew
rlabel  s 9 1 10 6 6 C0
port 1 nsew
rlabel  s 8 6 9 11 6 C0
port 1 nsew
rlabel  s 8 1 9 6 6 C0
port 1 nsew
rlabel  s 7 6 7 11 6 C0
port 1 nsew
rlabel  s 7 1 7 6 6 C0
port 1 nsew
rlabel  s 5 6 6 11 6 C0
port 1 nsew
rlabel  s 5 1 6 6 6 C0
port 1 nsew
rlabel  s 4 6 4 11 6 C0
port 1 nsew
rlabel  s 4 1 4 6 6 C0
port 1 nsew
rlabel  s 3 6 3 11 6 C0
port 1 nsew
rlabel  s 3 1 3 6 6 C0
port 1 nsew
rlabel  s 2 6 2 11 6 C0
port 1 nsew
rlabel  s 2 6 10 6 6 C0
port 1 nsew
rlabel  s 2 1 2 6 6 C0
port 1 nsew
rlabel  s 0 0 1 12 4 C0
port 1 nsew
rlabel  s 10 1 10 11 6 C1
port 2 nsew
rlabel  s 9 6 9 11 6 C1
port 2 nsew
rlabel  s 9 1 9 5 6 C1
port 2 nsew
rlabel  s 8 6 8 11 6 C1
port 2 nsew
rlabel  s 8 1 8 5 6 C1
port 2 nsew
rlabel  s 6 6 7 11 6 C1
port 2 nsew
rlabel  s 6 1 7 5 6 C1
port 2 nsew
rlabel  s 5 6 5 11 6 C1
port 2 nsew
rlabel  s 5 1 5 5 6 C1
port 2 nsew
rlabel  s 3 6 4 11 6 C1
port 2 nsew
rlabel  s 3 1 4 5 6 C1
port 2 nsew
rlabel  s 2 6 2 11 6 C1
port 2 nsew
rlabel  s 2 1 2 5 6 C1
port 2 nsew
rlabel  s 1 11 10 11 6 C1
port 2 nsew
rlabel  s 1 11 10 11 6 C1
port 2 nsew
rlabel  s 1 1 1 11 6 C1
port 2 nsew
rlabel  s 1 0 10 1 8 C1
port 2 nsew
rlabel r s 0 0 11 12 6 MET5
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 11 12
string LEFview TRUE
<< end >>
