magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s -3 -3 63 73 6 PAD
port 1 nsew
rlabel pfet_brown s -3 -3 63 -1 8 PAD
port 1 nsew
rlabel pfet_brown s 61 -1 63 71 6 PAD
port 1 nsew
rlabel pfet_brown s -3 -1 -1 71 4 PAD
port 1 nsew
rlabel pfet_brown s -3 71 63 73 6 PAD
port 1 nsew
rlabel  s -3 -3 63 0 8 PAD
port 1 nsew
rlabel  s 60 0 63 70 6 PAD
port 1 nsew
rlabel  s -3 0 0 70 4 PAD
port 1 nsew
rlabel  s -3 70 63 73 6 PAD
port 1 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -3 -3 62 72
string LEFview TRUE
<< end >>
