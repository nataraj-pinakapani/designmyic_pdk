magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel rotate s 2 6 2 6 6 GATE
port 1 nsew
rlabel rotate s 2 0 2 0 8 GATE
port 1 nsew
rlabel rotate s 1 6 1 6 6 GATE
port 1 nsew
rlabel rotate s 1 0 1 0 8 GATE
port 1 nsew
rlabel rotate s 1 6 1 6 6 GATE
port 1 nsew
rlabel rotate s 1 0 1 0 8 GATE
port 1 nsew
rlabel  s 1 6 2 6 6 GATE
port 2 nsew
rlabel  s 1 0 2 0 8 GATE
port 2 nsew
rlabel  s 1 6 2 6 6 GATE
port 2 nsew
rlabel  s 1 0 2 0 8 GATE
port 2 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 3 6
string LEFview TRUE
<< end >>
