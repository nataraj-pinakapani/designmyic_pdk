magic
tech minimum
timestamp 1644097873
<< properties >>
string gencell sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
string parameter m=1
string library sky130
<< end >>
