magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 4002 897
rect 3185 343 3698 377
<< pwell >>
rect 1545 283 1967 290
rect 1041 217 1967 283
rect 2408 217 3435 283
rect 3666 217 3932 283
rect 86 43 3932 217
rect -26 -43 3962 43
<< mvnmos >>
rect 169 107 269 191
rect 325 107 425 191
rect 467 107 567 191
rect 623 107 723 191
rect 765 107 865 191
rect 1124 107 1224 257
rect 1354 173 1454 257
rect 1628 180 1728 264
rect 1784 180 1884 264
rect 2058 107 2158 191
rect 2214 107 2314 191
rect 2491 173 2591 257
rect 2647 173 2747 257
rect 2789 173 2889 257
rect 2968 107 3068 257
rect 3252 107 3352 257
rect 3431 107 3531 191
rect 3749 107 3849 257
<< mvpmos >>
rect 325 659 425 743
rect 481 659 581 743
rect 83 515 183 599
rect 747 598 847 682
rect 903 598 1003 682
rect 1169 543 1269 743
rect 1428 579 1528 663
rect 1570 579 1670 663
rect 1726 579 1826 663
rect 1996 468 2096 618
rect 2152 468 2252 618
rect 2418 445 2518 529
rect 2593 445 2693 645
rect 2863 543 2963 627
rect 3038 543 3138 743
rect 3304 409 3404 709
rect 3479 409 3579 559
rect 3749 443 3849 743
<< mvndiff >>
rect 1067 249 1124 257
rect 1067 215 1079 249
rect 1113 215 1124 249
rect 112 166 169 191
rect 112 132 124 166
rect 158 132 169 166
rect 112 107 169 132
rect 269 166 325 191
rect 269 132 280 166
rect 314 132 325 166
rect 269 107 325 132
rect 425 107 467 191
rect 567 166 623 191
rect 567 132 578 166
rect 612 132 623 166
rect 567 107 623 132
rect 723 107 765 191
rect 865 166 922 191
rect 865 132 876 166
rect 910 132 922 166
rect 865 107 922 132
rect 1067 157 1124 215
rect 1067 123 1079 157
rect 1113 123 1124 157
rect 1067 107 1124 123
rect 1224 182 1354 257
rect 1224 148 1251 182
rect 1285 173 1354 182
rect 1454 215 1511 257
rect 1454 181 1465 215
rect 1499 181 1511 215
rect 1454 173 1511 181
rect 1571 239 1628 264
rect 1571 205 1583 239
rect 1617 205 1628 239
rect 1571 180 1628 205
rect 1728 239 1784 264
rect 1728 205 1739 239
rect 1773 205 1784 239
rect 1728 180 1784 205
rect 1884 239 1941 264
rect 1884 205 1895 239
rect 1929 205 1941 239
rect 1884 180 1941 205
rect 2434 232 2491 257
rect 2434 198 2446 232
rect 2480 198 2491 232
rect 1285 148 1297 173
rect 1224 107 1297 148
rect 2001 166 2058 191
rect 2001 132 2013 166
rect 2047 132 2058 166
rect 2001 107 2058 132
rect 2158 166 2214 191
rect 2158 132 2169 166
rect 2203 132 2214 166
rect 2158 107 2214 132
rect 2314 166 2371 191
rect 2434 173 2491 198
rect 2591 232 2647 257
rect 2591 198 2602 232
rect 2636 198 2647 232
rect 2591 173 2647 198
rect 2747 173 2789 257
rect 2889 249 2968 257
rect 2889 215 2923 249
rect 2957 215 2968 249
rect 2889 173 2968 215
rect 2314 132 2325 166
rect 2359 132 2371 166
rect 2911 149 2968 173
rect 2314 107 2371 132
rect 2911 115 2923 149
rect 2957 115 2968 149
rect 2911 107 2968 115
rect 3068 249 3125 257
rect 3068 215 3079 249
rect 3113 215 3125 249
rect 3068 149 3125 215
rect 3068 115 3079 149
rect 3113 115 3125 149
rect 3068 107 3125 115
rect 3195 249 3252 257
rect 3195 215 3207 249
rect 3241 215 3252 249
rect 3195 149 3252 215
rect 3195 115 3207 149
rect 3241 115 3252 149
rect 3195 107 3252 115
rect 3352 249 3409 257
rect 3352 215 3363 249
rect 3397 215 3409 249
rect 3352 191 3409 215
rect 3692 249 3749 257
rect 3692 215 3704 249
rect 3738 215 3749 249
rect 3352 149 3431 191
rect 3352 115 3363 149
rect 3397 115 3431 149
rect 3352 107 3431 115
rect 3531 166 3588 191
rect 3531 132 3542 166
rect 3576 132 3588 166
rect 3531 107 3588 132
rect 3692 149 3749 215
rect 3692 115 3704 149
rect 3738 115 3749 149
rect 3692 107 3749 115
rect 3849 249 3906 257
rect 3849 215 3860 249
rect 3894 215 3906 249
rect 3849 149 3906 215
rect 3849 115 3860 149
rect 3894 115 3906 149
rect 3849 107 3906 115
<< mvpdiff >>
rect 268 718 325 743
rect 268 684 280 718
rect 314 684 325 718
rect 268 659 325 684
rect 425 718 481 743
rect 425 684 436 718
rect 470 684 481 718
rect 425 659 481 684
rect 581 718 634 743
rect 581 684 592 718
rect 626 684 634 718
rect 581 659 634 684
rect 30 574 83 599
rect 30 540 38 574
rect 72 540 83 574
rect 30 515 83 540
rect 183 574 240 599
rect 183 540 194 574
rect 228 540 240 574
rect 183 515 240 540
rect 694 657 747 682
rect 694 623 702 657
rect 736 623 747 657
rect 694 598 747 623
rect 847 657 903 682
rect 847 623 858 657
rect 892 623 903 657
rect 847 598 903 623
rect 1003 657 1056 682
rect 1003 623 1014 657
rect 1048 623 1056 657
rect 1003 598 1056 623
rect 1116 675 1169 743
rect 1116 641 1124 675
rect 1158 641 1169 675
rect 1116 589 1169 641
rect 1116 555 1124 589
rect 1158 555 1169 589
rect 1116 543 1169 555
rect 1269 731 1326 743
rect 1269 697 1280 731
rect 1314 697 1326 731
rect 1269 663 1326 697
rect 2985 731 3038 743
rect 2985 697 2993 731
rect 3027 697 3038 731
rect 1269 579 1428 663
rect 1528 579 1570 663
rect 1670 621 1726 663
rect 1670 587 1681 621
rect 1715 587 1726 621
rect 1670 579 1726 587
rect 1826 654 1883 663
rect 1826 620 1837 654
rect 1871 620 1883 654
rect 2985 660 3038 697
rect 1826 579 1883 620
rect 2540 621 2593 645
rect 1269 543 1326 579
rect 1943 514 1996 618
rect 1943 480 1951 514
rect 1985 480 1996 514
rect 1943 468 1996 480
rect 2096 595 2152 618
rect 2096 561 2107 595
rect 2141 561 2152 595
rect 2096 468 2152 561
rect 2252 606 2305 618
rect 2252 572 2263 606
rect 2297 572 2305 606
rect 2252 514 2305 572
rect 2540 587 2548 621
rect 2582 587 2593 621
rect 2540 529 2593 587
rect 2252 480 2263 514
rect 2297 480 2305 514
rect 2252 468 2305 480
rect 2365 504 2418 529
rect 2365 470 2373 504
rect 2407 470 2418 504
rect 2365 445 2418 470
rect 2518 491 2593 529
rect 2518 457 2548 491
rect 2582 457 2593 491
rect 2518 445 2593 457
rect 2693 637 2750 645
rect 2693 603 2704 637
rect 2738 603 2750 637
rect 2985 627 2993 660
rect 2693 562 2750 603
rect 2693 528 2704 562
rect 2738 528 2750 562
rect 2810 602 2863 627
rect 2810 568 2818 602
rect 2852 568 2863 602
rect 2810 543 2863 568
rect 2963 626 2993 627
rect 3027 626 3038 660
rect 2963 589 3038 626
rect 2963 555 2993 589
rect 3027 555 3038 589
rect 2963 543 3038 555
rect 3138 731 3191 743
rect 3692 735 3749 743
rect 3138 697 3149 731
rect 3183 697 3191 731
rect 3138 660 3191 697
rect 3138 626 3149 660
rect 3183 626 3191 660
rect 3138 589 3191 626
rect 3138 555 3149 589
rect 3183 555 3191 589
rect 3138 543 3191 555
rect 3251 691 3304 709
rect 3251 657 3259 691
rect 3293 657 3304 691
rect 3251 613 3304 657
rect 3251 579 3259 613
rect 3293 579 3304 613
rect 2693 487 2750 528
rect 2693 453 2704 487
rect 2738 453 2750 487
rect 2693 445 2750 453
rect 3251 533 3304 579
rect 3251 499 3259 533
rect 3293 499 3304 533
rect 3251 455 3304 499
rect 3251 421 3259 455
rect 3293 421 3304 455
rect 3251 409 3304 421
rect 3404 697 3457 709
rect 3404 663 3415 697
rect 3449 663 3457 697
rect 3404 617 3457 663
rect 3404 583 3415 617
rect 3449 583 3457 617
rect 3692 701 3704 735
rect 3738 701 3749 735
rect 3692 652 3749 701
rect 3692 618 3704 652
rect 3738 618 3749 652
rect 3404 559 3457 583
rect 3692 568 3749 618
rect 3404 535 3479 559
rect 3404 501 3415 535
rect 3449 501 3479 535
rect 3404 455 3479 501
rect 3404 421 3415 455
rect 3449 421 3479 455
rect 3404 409 3479 421
rect 3579 547 3632 559
rect 3579 513 3590 547
rect 3624 513 3632 547
rect 3579 455 3632 513
rect 3579 421 3590 455
rect 3624 421 3632 455
rect 3692 534 3704 568
rect 3738 534 3749 568
rect 3692 485 3749 534
rect 3692 451 3704 485
rect 3738 451 3749 485
rect 3692 443 3749 451
rect 3849 735 3906 743
rect 3849 701 3860 735
rect 3894 701 3906 735
rect 3849 652 3906 701
rect 3849 618 3860 652
rect 3894 618 3906 652
rect 3849 568 3906 618
rect 3849 534 3860 568
rect 3894 534 3906 568
rect 3849 485 3906 534
rect 3849 451 3860 485
rect 3894 451 3906 485
rect 3849 443 3906 451
rect 3579 409 3632 421
<< mvndiffc >>
rect 1079 215 1113 249
rect 124 132 158 166
rect 280 132 314 166
rect 578 132 612 166
rect 876 132 910 166
rect 1079 123 1113 157
rect 1251 148 1285 182
rect 1465 181 1499 215
rect 1583 205 1617 239
rect 1739 205 1773 239
rect 1895 205 1929 239
rect 2446 198 2480 232
rect 2013 132 2047 166
rect 2169 132 2203 166
rect 2602 198 2636 232
rect 2923 215 2957 249
rect 2325 132 2359 166
rect 2923 115 2957 149
rect 3079 215 3113 249
rect 3079 115 3113 149
rect 3207 215 3241 249
rect 3207 115 3241 149
rect 3363 215 3397 249
rect 3704 215 3738 249
rect 3363 115 3397 149
rect 3542 132 3576 166
rect 3704 115 3738 149
rect 3860 215 3894 249
rect 3860 115 3894 149
<< mvpdiffc >>
rect 280 684 314 718
rect 436 684 470 718
rect 592 684 626 718
rect 38 540 72 574
rect 194 540 228 574
rect 702 623 736 657
rect 858 623 892 657
rect 1014 623 1048 657
rect 1124 641 1158 675
rect 1124 555 1158 589
rect 1280 697 1314 731
rect 2993 697 3027 731
rect 1681 587 1715 621
rect 1837 620 1871 654
rect 1951 480 1985 514
rect 2107 561 2141 595
rect 2263 572 2297 606
rect 2548 587 2582 621
rect 2263 480 2297 514
rect 2373 470 2407 504
rect 2548 457 2582 491
rect 2704 603 2738 637
rect 2704 528 2738 562
rect 2818 568 2852 602
rect 2993 626 3027 660
rect 2993 555 3027 589
rect 3149 697 3183 731
rect 3149 626 3183 660
rect 3149 555 3183 589
rect 3259 657 3293 691
rect 3259 579 3293 613
rect 2704 453 2738 487
rect 3259 499 3293 533
rect 3259 421 3293 455
rect 3415 663 3449 697
rect 3415 583 3449 617
rect 3704 701 3738 735
rect 3704 618 3738 652
rect 3415 501 3449 535
rect 3415 421 3449 455
rect 3590 513 3624 547
rect 3590 421 3624 455
rect 3704 534 3738 568
rect 3704 451 3738 485
rect 3860 701 3894 735
rect 3860 618 3894 652
rect 3860 534 3894 568
rect 3860 451 3894 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3936 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3936 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
<< poly >>
rect 325 743 425 769
rect 481 743 581 769
rect 1169 743 1269 769
rect 3038 743 3138 769
rect 3749 743 3849 769
rect 747 682 847 708
rect 903 682 1003 708
rect 83 599 183 625
rect 83 448 183 515
rect 325 488 425 659
rect 481 557 581 659
rect 747 572 847 598
rect 325 454 345 488
rect 379 454 425 488
rect 83 428 269 448
rect 83 394 129 428
rect 163 394 269 428
rect 83 360 269 394
rect 83 326 129 360
rect 163 326 269 360
rect 83 217 269 326
rect 169 191 269 217
rect 325 420 425 454
rect 325 386 345 420
rect 379 386 425 420
rect 325 191 425 386
rect 467 537 581 557
rect 467 503 501 537
rect 535 503 581 537
rect 467 469 581 503
rect 467 435 501 469
rect 535 435 581 469
rect 467 415 581 435
rect 623 472 847 572
rect 467 191 567 415
rect 623 373 723 472
rect 903 373 1003 598
rect 1428 663 1528 689
rect 1570 663 1670 689
rect 1726 663 1826 689
rect 2593 645 2693 671
rect 1996 618 2096 644
rect 2152 618 2252 644
rect 1169 521 1269 543
rect 609 353 723 373
rect 609 319 629 353
rect 663 319 723 353
rect 609 285 723 319
rect 609 251 629 285
rect 663 251 723 285
rect 609 217 723 251
rect 623 191 723 217
rect 765 353 1003 373
rect 765 319 849 353
rect 883 319 1003 353
rect 765 285 1003 319
rect 765 251 849 285
rect 883 251 1003 285
rect 1124 495 1334 521
rect 1124 461 1280 495
rect 1314 461 1334 495
rect 1124 421 1334 461
rect 1124 279 1269 421
rect 1428 379 1528 579
rect 1570 557 1670 579
rect 1570 531 1684 557
rect 1570 497 1634 531
rect 1668 497 1684 531
rect 1570 457 1684 497
rect 1354 355 1528 379
rect 1354 321 1374 355
rect 1408 321 1528 355
rect 1354 279 1528 321
rect 1584 386 1684 457
rect 1726 553 1826 579
rect 1726 453 1884 553
rect 2418 529 2518 555
rect 1784 427 1884 453
rect 1784 393 1830 427
rect 1864 393 1884 427
rect 1584 286 1728 386
rect 1124 257 1224 279
rect 1354 257 1454 279
rect 1628 264 1728 286
rect 1784 359 1884 393
rect 1784 325 1830 359
rect 1864 325 1884 359
rect 1784 264 1884 325
rect 1996 420 2096 468
rect 1996 386 2021 420
rect 2055 386 2096 420
rect 1996 309 2096 386
rect 2152 446 2252 468
rect 2152 419 2314 446
rect 2863 627 2963 653
rect 3304 709 3404 735
rect 2863 521 2963 543
rect 2789 495 2963 521
rect 2789 461 2909 495
rect 2943 461 2963 495
rect 2418 419 2518 445
rect 2152 385 2172 419
rect 2206 385 2314 419
rect 2152 351 2314 385
rect 1996 267 2169 309
rect 765 217 1003 251
rect 765 191 865 217
rect 1996 233 2115 267
rect 2149 233 2169 267
rect 1996 213 2169 233
rect 2058 191 2158 213
rect 2214 191 2314 351
rect 2356 397 2518 419
rect 2356 363 2376 397
rect 2410 363 2518 397
rect 2593 423 2693 445
rect 2593 379 2739 423
rect 2789 421 2963 461
rect 2593 372 2747 379
rect 2356 330 2518 363
rect 2639 341 2747 372
rect 2356 329 2591 330
rect 2356 295 2376 329
rect 2410 295 2591 329
rect 2356 279 2591 295
rect 2639 307 2672 341
rect 2706 307 2747 341
rect 2639 279 2747 307
rect 2491 257 2591 279
rect 2647 257 2747 279
rect 2789 257 2889 421
rect 3038 379 3138 543
rect 3479 559 3579 585
rect 3749 417 3849 443
rect 3304 383 3404 409
rect 3479 383 3579 409
rect 2957 359 3138 379
rect 2957 325 2977 359
rect 3011 325 3138 359
rect 2957 279 3138 325
rect 3252 351 3579 383
rect 3252 317 3361 351
rect 3395 317 3579 351
rect 3252 283 3579 317
rect 3738 351 3849 417
rect 3738 317 3758 351
rect 3792 317 3849 351
rect 3738 283 3849 317
rect 2968 257 3068 279
rect 3252 257 3352 283
rect 1354 147 1454 173
rect 1628 154 1728 180
rect 1784 154 1884 180
rect 2491 147 2591 173
rect 2647 147 2747 173
rect 2789 147 2889 173
rect 3431 191 3531 283
rect 3749 257 3849 283
rect 169 81 269 107
rect 325 81 425 107
rect 467 81 567 107
rect 623 81 723 107
rect 765 81 865 107
rect 1124 81 1224 107
rect 2058 81 2158 107
rect 2214 81 2314 107
rect 2968 81 3068 107
rect 3252 81 3352 107
rect 3431 81 3531 107
rect 3749 81 3849 107
<< polycont >>
rect 345 454 379 488
rect 129 394 163 428
rect 129 326 163 360
rect 345 386 379 420
rect 501 503 535 537
rect 501 435 535 469
rect 629 319 663 353
rect 629 251 663 285
rect 849 319 883 353
rect 849 251 883 285
rect 1280 461 1314 495
rect 1634 497 1668 531
rect 1374 321 1408 355
rect 1830 393 1864 427
rect 1830 325 1864 359
rect 2021 386 2055 420
rect 2909 461 2943 495
rect 2172 385 2206 419
rect 2115 233 2149 267
rect 2376 363 2410 397
rect 2376 295 2410 329
rect 2672 307 2706 341
rect 2977 325 3011 359
rect 3361 317 3395 351
rect 3758 317 3792 351
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3936 831
rect 126 735 244 741
rect 126 701 132 735
rect 166 701 204 735
rect 238 701 244 735
rect 22 574 88 603
rect 22 540 38 574
rect 72 540 88 574
rect 22 511 88 540
rect 126 574 244 701
rect 280 718 314 751
rect 280 619 314 684
rect 350 735 540 751
rect 350 701 356 735
rect 390 701 428 735
rect 462 718 500 735
rect 470 701 500 718
rect 534 701 540 735
rect 350 684 436 701
rect 470 684 540 701
rect 350 667 540 684
rect 576 722 806 756
rect 576 718 642 722
rect 576 684 592 718
rect 626 684 642 718
rect 576 655 642 684
rect 686 657 736 686
rect 686 623 702 657
rect 686 619 736 623
rect 280 585 736 619
rect 126 540 194 574
rect 228 540 244 574
rect 772 570 806 722
rect 842 727 1228 761
rect 842 657 908 727
rect 842 623 858 657
rect 892 623 908 657
rect 842 606 908 623
rect 998 657 1048 686
rect 998 623 1014 657
rect 998 570 1048 623
rect 126 524 244 540
rect 485 537 551 549
rect 22 269 56 511
rect 485 503 501 537
rect 535 503 551 537
rect 772 536 1048 570
rect 1084 675 1158 691
rect 1084 646 1124 675
rect 1084 612 1087 646
rect 1121 641 1124 646
rect 1121 612 1158 641
rect 1084 589 1158 612
rect 1084 555 1124 589
rect 313 454 345 488
rect 379 454 395 488
rect 113 428 179 444
rect 113 394 129 428
rect 163 394 179 428
rect 113 360 179 394
rect 313 420 395 454
rect 313 386 345 420
rect 379 386 395 420
rect 485 469 551 503
rect 485 435 501 469
rect 535 435 551 469
rect 113 326 129 360
rect 163 350 179 360
rect 485 350 551 435
rect 702 466 1027 500
rect 163 326 551 350
rect 113 310 551 326
rect 613 353 666 369
rect 613 319 629 353
rect 663 319 666 353
rect 613 285 666 319
rect 613 269 629 285
rect 22 251 629 269
rect 663 251 666 285
rect 22 235 666 251
rect 108 166 174 235
rect 702 199 736 466
rect 833 353 935 430
rect 833 319 849 353
rect 883 319 935 353
rect 833 285 935 319
rect 833 251 849 285
rect 883 251 935 285
rect 833 235 935 251
rect 108 132 124 166
rect 158 132 174 166
rect 108 99 174 132
rect 210 166 400 199
rect 210 132 280 166
rect 314 132 400 166
rect 210 113 400 132
rect 210 79 216 113
rect 250 79 288 113
rect 322 79 360 113
rect 394 79 400 113
rect 562 166 736 199
rect 562 132 578 166
rect 612 165 736 166
rect 772 166 957 199
rect 612 132 628 165
rect 562 99 628 132
rect 772 132 876 166
rect 910 132 957 166
rect 772 113 957 132
rect 210 73 400 79
rect 772 79 775 113
rect 809 79 847 113
rect 881 79 919 113
rect 953 79 957 113
rect 772 73 957 79
rect 993 87 1027 466
rect 1084 355 1158 555
rect 1194 657 1228 727
rect 1264 735 1442 751
rect 1298 731 1336 735
rect 1314 701 1336 731
rect 1370 701 1408 735
rect 1264 697 1280 701
rect 1314 697 1442 701
rect 1264 693 1442 697
rect 2107 735 2225 741
rect 2107 701 2113 735
rect 2147 701 2185 735
rect 2219 701 2225 735
rect 1478 657 1887 691
rect 1194 623 1512 657
rect 1821 654 1887 657
rect 1194 425 1228 623
rect 1548 587 1681 621
rect 1715 587 1731 621
rect 1821 620 1837 654
rect 1871 620 1887 654
rect 1548 571 1731 587
rect 2107 595 2225 701
rect 2357 727 2868 761
rect 1548 511 1582 571
rect 1767 550 2071 584
rect 1767 535 1801 550
rect 1264 495 1582 511
rect 1618 531 1801 535
rect 1618 497 1634 531
rect 1668 497 1801 531
rect 1264 461 1280 495
rect 1314 461 1582 495
rect 1935 480 1951 514
rect 1985 480 2001 514
rect 1935 464 2001 480
rect 2037 494 2071 550
rect 2141 561 2225 595
rect 2107 530 2225 561
rect 2263 606 2313 622
rect 2297 572 2313 606
rect 2263 514 2313 572
rect 2037 480 2263 494
rect 2297 480 2313 514
rect 1548 427 1757 461
rect 1194 391 1494 425
rect 1063 321 1374 355
rect 1408 321 1424 355
rect 1063 249 1129 321
rect 1460 285 1494 391
rect 1063 215 1079 249
rect 1113 215 1129 249
rect 1063 157 1129 215
rect 1063 123 1079 157
rect 1113 123 1129 157
rect 1165 251 1633 285
rect 1165 87 1199 251
rect 1567 239 1633 251
rect 993 53 1199 87
rect 1235 182 1413 215
rect 1235 148 1251 182
rect 1285 148 1413 182
rect 1235 113 1413 148
rect 1449 181 1465 215
rect 1499 181 1515 215
rect 1567 205 1583 239
rect 1617 205 1633 239
rect 1567 188 1633 205
rect 1723 272 1757 427
rect 1814 427 1880 443
rect 1814 393 1830 427
rect 1864 393 1880 427
rect 1814 359 1880 393
rect 1814 325 1830 359
rect 1864 343 1880 359
rect 1935 343 1969 464
rect 2037 460 2313 480
rect 2357 504 2423 727
rect 2357 470 2373 504
rect 2407 470 2423 504
rect 2037 428 2071 460
rect 2357 441 2423 470
rect 2462 657 2759 691
rect 2005 420 2071 428
rect 2005 386 2021 420
rect 2055 386 2071 420
rect 2005 379 2071 386
rect 2137 419 2279 424
rect 2137 385 2172 419
rect 2206 385 2279 419
rect 2137 379 2279 385
rect 2360 397 2426 405
rect 2360 363 2376 397
rect 2410 363 2426 397
rect 2360 343 2426 363
rect 1864 329 2426 343
rect 1864 325 2376 329
rect 1814 309 2376 325
rect 1723 239 1789 272
rect 1723 205 1739 239
rect 1773 205 1789 239
rect 1723 188 1789 205
rect 1879 239 1945 272
rect 1879 205 1895 239
rect 1929 205 1945 239
rect 1449 152 1515 181
rect 1879 152 1945 205
rect 1449 118 1945 152
rect 1997 166 2063 309
rect 2360 295 2376 309
rect 2410 295 2426 329
rect 2360 289 2426 295
rect 2099 267 2165 273
rect 2099 233 2115 267
rect 2149 253 2165 267
rect 2149 233 2375 253
rect 2462 249 2496 657
rect 2688 646 2759 657
rect 2688 637 2719 646
rect 2532 587 2548 621
rect 2582 587 2598 621
rect 2532 491 2598 587
rect 2532 457 2548 491
rect 2582 457 2598 491
rect 2532 441 2598 457
rect 2688 603 2704 637
rect 2753 612 2759 646
rect 2738 603 2759 612
rect 2688 562 2759 603
rect 2688 528 2704 562
rect 2738 528 2759 562
rect 2802 602 2868 727
rect 2802 568 2818 602
rect 2852 568 2868 602
rect 2802 539 2868 568
rect 2904 735 3085 747
rect 2904 701 2905 735
rect 2939 701 2977 735
rect 3011 731 3049 735
rect 3027 701 3049 731
rect 3083 701 3085 735
rect 2904 697 2993 701
rect 3027 697 3085 701
rect 2904 660 3085 697
rect 2904 626 2993 660
rect 3027 626 3085 660
rect 2904 589 3085 626
rect 2904 555 2993 589
rect 3027 555 3085 589
rect 2904 539 3085 555
rect 3121 731 3379 761
rect 3121 697 3149 731
rect 3183 727 3379 731
rect 3183 697 3199 727
rect 3121 660 3199 697
rect 3121 626 3149 660
rect 3183 626 3199 660
rect 3121 589 3199 626
rect 3121 555 3149 589
rect 3183 555 3199 589
rect 3121 539 3199 555
rect 3243 657 3259 691
rect 3293 657 3309 691
rect 3243 613 3309 657
rect 3243 579 3259 613
rect 3293 579 3309 613
rect 2688 487 2759 528
rect 3121 503 3155 539
rect 3243 533 3309 579
rect 3243 503 3259 533
rect 2688 453 2704 487
rect 2738 453 2759 487
rect 2893 495 3155 503
rect 2893 461 2909 495
rect 2943 461 3155 495
rect 2893 453 3155 461
rect 2099 219 2375 233
rect 1997 132 2013 166
rect 2047 132 2063 166
rect 1269 79 1307 113
rect 1341 79 1379 113
rect 1997 99 2063 132
rect 2099 166 2289 183
rect 2099 132 2169 166
rect 2203 132 2289 166
rect 2099 113 2289 132
rect 1235 73 1413 79
rect 2099 79 2105 113
rect 2139 79 2177 113
rect 2211 79 2249 113
rect 2283 79 2289 113
rect 2325 166 2375 219
rect 2359 132 2375 166
rect 2430 232 2496 249
rect 2430 198 2446 232
rect 2480 198 2496 232
rect 2430 165 2496 198
rect 2564 417 2598 441
rect 2564 383 3027 417
rect 2564 265 2598 383
rect 2961 359 3027 383
rect 2656 341 2722 347
rect 2656 307 2672 341
rect 2706 307 2722 341
rect 2961 325 2977 359
rect 3011 325 3027 359
rect 2961 309 3027 325
rect 2656 301 2722 307
rect 2564 232 2652 265
rect 2564 198 2602 232
rect 2636 198 2652 232
rect 2564 165 2652 198
rect 2325 129 2375 132
rect 2688 129 2722 301
rect 2325 95 2722 129
rect 2783 249 2973 265
rect 2783 215 2923 249
rect 2957 215 2973 249
rect 2783 149 2973 215
rect 2783 115 2923 149
rect 2957 115 2973 149
rect 2783 113 2973 115
rect 2099 73 2289 79
rect 2783 79 2789 113
rect 2823 79 2861 113
rect 2895 79 2933 113
rect 2967 79 2973 113
rect 3063 249 3155 453
rect 3063 215 3079 249
rect 3113 215 3155 249
rect 3063 149 3155 215
rect 3063 115 3079 149
rect 3113 115 3155 149
rect 3063 99 3155 115
rect 3191 499 3259 503
rect 3293 499 3309 533
rect 3191 455 3309 499
rect 3191 421 3259 455
rect 3293 421 3309 455
rect 3191 405 3309 421
rect 3191 249 3257 405
rect 3345 367 3379 727
rect 3415 735 3533 741
rect 3415 701 3421 735
rect 3455 701 3493 735
rect 3527 701 3533 735
rect 3415 697 3533 701
rect 3449 663 3533 697
rect 3415 617 3533 663
rect 3449 583 3533 617
rect 3415 535 3533 583
rect 3676 735 3794 751
rect 3676 701 3682 735
rect 3738 701 3754 735
rect 3788 701 3794 735
rect 3676 652 3794 701
rect 3676 618 3704 652
rect 3738 618 3794 652
rect 3676 568 3794 618
rect 3449 501 3533 535
rect 3415 455 3533 501
rect 3449 421 3533 455
rect 3415 405 3533 421
rect 3574 547 3640 563
rect 3574 513 3590 547
rect 3624 513 3640 547
rect 3574 455 3640 513
rect 3574 421 3590 455
rect 3624 421 3640 455
rect 3676 534 3704 568
rect 3738 534 3794 568
rect 3676 485 3794 534
rect 3676 451 3704 485
rect 3738 451 3794 485
rect 3676 435 3794 451
rect 3844 735 3911 751
rect 3844 701 3860 735
rect 3894 701 3911 735
rect 3844 652 3911 701
rect 3844 618 3860 652
rect 3894 618 3911 652
rect 3844 568 3911 618
rect 3844 534 3860 568
rect 3894 534 3911 568
rect 3844 485 3911 534
rect 3844 451 3860 485
rect 3894 451 3911 485
rect 3574 405 3640 421
rect 3606 367 3640 405
rect 3345 351 3411 367
rect 3345 317 3361 351
rect 3395 317 3411 351
rect 3606 351 3808 367
rect 3606 335 3758 351
rect 3345 301 3411 317
rect 3526 317 3758 335
rect 3792 317 3808 351
rect 3526 301 3808 317
rect 3191 215 3207 249
rect 3241 215 3257 249
rect 3191 149 3257 215
rect 3191 115 3207 149
rect 3241 115 3257 149
rect 3191 99 3257 115
rect 3293 249 3483 265
rect 3293 215 3363 249
rect 3397 215 3483 249
rect 3293 149 3483 215
rect 3293 115 3363 149
rect 3397 115 3483 149
rect 3293 113 3483 115
rect 2783 73 2973 79
rect 3293 79 3299 113
rect 3333 79 3371 113
rect 3405 79 3443 113
rect 3477 79 3483 113
rect 3526 166 3592 301
rect 3526 132 3542 166
rect 3576 132 3592 166
rect 3526 99 3592 132
rect 3628 249 3808 265
rect 3628 215 3704 249
rect 3738 215 3808 249
rect 3628 149 3808 215
rect 3628 115 3704 149
rect 3738 115 3808 149
rect 3628 113 3808 115
rect 3293 73 3483 79
rect 3628 79 3629 113
rect 3663 79 3701 113
rect 3735 79 3773 113
rect 3807 79 3808 113
rect 3844 249 3911 451
rect 3844 215 3860 249
rect 3894 215 3911 249
rect 3844 149 3911 215
rect 3844 115 3860 149
rect 3894 115 3911 149
rect 3844 99 3911 115
rect 3628 73 3808 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3936 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 132 701 166 735
rect 204 701 238 735
rect 356 701 390 735
rect 428 718 462 735
rect 428 701 436 718
rect 436 701 462 718
rect 500 701 534 735
rect 1087 612 1121 646
rect 216 79 250 113
rect 288 79 322 113
rect 360 79 394 113
rect 775 79 809 113
rect 847 79 881 113
rect 919 79 953 113
rect 1264 731 1298 735
rect 1264 701 1280 731
rect 1280 701 1298 731
rect 1336 701 1370 735
rect 1408 701 1442 735
rect 2113 701 2147 735
rect 2185 701 2219 735
rect 2719 637 2753 646
rect 2719 612 2738 637
rect 2738 612 2753 637
rect 2905 701 2939 735
rect 2977 731 3011 735
rect 2977 701 2993 731
rect 2993 701 3011 731
rect 3049 701 3083 735
rect 1235 79 1269 113
rect 1307 79 1341 113
rect 1379 79 1413 113
rect 2105 79 2139 113
rect 2177 79 2211 113
rect 2249 79 2283 113
rect 2789 79 2823 113
rect 2861 79 2895 113
rect 2933 79 2967 113
rect 3421 701 3455 735
rect 3493 701 3527 735
rect 3682 701 3704 735
rect 3704 701 3716 735
rect 3754 701 3788 735
rect 3299 79 3333 113
rect 3371 79 3405 113
rect 3443 79 3477 113
rect 3629 79 3663 113
rect 3701 79 3735 113
rect 3773 79 3807 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
<< metal1 >>
rect 0 831 3936 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3936 831
rect 0 791 3936 797
rect 0 735 3936 763
rect 0 701 132 735
rect 166 701 204 735
rect 238 701 356 735
rect 390 701 428 735
rect 462 701 500 735
rect 534 701 1264 735
rect 1298 701 1336 735
rect 1370 701 1408 735
rect 1442 701 2113 735
rect 2147 701 2185 735
rect 2219 701 2905 735
rect 2939 701 2977 735
rect 3011 701 3049 735
rect 3083 701 3421 735
rect 3455 701 3493 735
rect 3527 701 3682 735
rect 3716 701 3754 735
rect 3788 701 3936 735
rect 0 689 3936 701
rect 1075 646 1133 652
rect 1075 612 1087 646
rect 1121 643 1133 646
rect 2707 646 2765 652
rect 2707 643 2719 646
rect 1121 615 2719 643
rect 1121 612 1133 615
rect 1075 606 1133 612
rect 2707 612 2719 615
rect 2753 612 2765 646
rect 2707 606 2765 612
rect 0 113 3936 125
rect 0 79 216 113
rect 250 79 288 113
rect 322 79 360 113
rect 394 79 775 113
rect 809 79 847 113
rect 881 79 919 113
rect 953 79 1235 113
rect 1269 79 1307 113
rect 1341 79 1379 113
rect 1413 79 2105 113
rect 2139 79 2177 113
rect 2211 79 2249 113
rect 2283 79 2789 113
rect 2823 79 2861 113
rect 2895 79 2933 113
rect 2967 79 3299 113
rect 3333 79 3371 113
rect 3405 79 3443 113
rect 3477 79 3629 113
rect 3663 79 3701 113
rect 3735 79 3773 113
rect 3807 79 3936 113
rect 0 51 3936 79
rect 0 17 3936 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3936 17
rect 0 -23 3936 -17
<< labels >>
flabel comment s 2055 332 2055 332 0 FreeSans 200 90 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfxbp_1
flabel metal1 s 0 51 3936 125 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 0 3936 23 0 FreeSans 340 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 0 689 3936 763 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 791 3936 814 0 FreeSans 340 0 0 0 VPB
port 7 nsew power bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3199 168 3233 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 3199 242 3233 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 3199 316 3233 350 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 3199 390 3233 424 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 3199 464 3233 498 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 3871 168 3905 202 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3871 242 3905 276 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3871 316 3905 350 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3871 390 3905 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3871 464 3905 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3871 538 3905 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3871 612 3905 646 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3936 814
string GDS_END 643078
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 605408
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
