magic
tech sky130B
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__hvdfm1sd2__example_5595914180827  sky130_fd_pr__hvdfm1sd2__example_5595914180827_0
timestamp 1663361622
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808233  sky130_fd_pr__hvdfm1sd__example_55959141808233_0
timestamp 1663361622
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808233  sky130_fd_pr__hvdfm1sd__example_55959141808233_1
timestamp 1663361622
transform 1 0 256 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 32670196
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 32668754
<< end >>
