/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/sky130_fd_pr__pfet_01v8_lvt_fail.cdl