magic
tech sky130B
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_0
timestamp 1663361622
transform -1 0 -80 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_1
timestamp 1663361622
transform 1 0 117 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 8136902
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 8135912
<< end >>
