magic
tech sky130A
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_0
timestamp 1663361622
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_1
timestamp 1663361622
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_2
timestamp 1663361622
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_3
timestamp 1663361622
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_4
timestamp 1663361622
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_5
timestamp 1663361622
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_6
timestamp 1663361622
transform 1 0 1036 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_7
timestamp 1663361622
transform 1 0 1192 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_8
timestamp 1663361622
transform 1 0 1348 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_9
timestamp 1663361622
transform 1 0 1504 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_10
timestamp 1663361622
transform 1 0 1660 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_11
timestamp 1663361622
transform 1 0 1816 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_12
timestamp 1663361622
transform 1 0 1972 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_13
timestamp 1663361622
transform 1 0 2128 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_14
timestamp 1663361622
transform 1 0 2284 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_15
timestamp 1663361622
transform 1 0 2440 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_16
timestamp 1663361622
transform 1 0 2596 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_17
timestamp 1663361622
transform 1 0 2752 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_18
timestamp 1663361622
transform 1 0 2908 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_19
timestamp 1663361622
transform 1 0 3064 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_20
timestamp 1663361622
transform 1 0 3220 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_21
timestamp 1663361622
transform 1 0 3376 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_22
timestamp 1663361622
transform 1 0 3532 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_23
timestamp 1663361622
transform 1 0 3688 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_24
timestamp 1663361622
transform 1 0 3844 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_25
timestamp 1663361622
transform 1 0 4000 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_26
timestamp 1663361622
transform 1 0 4156 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_27
timestamp 1663361622
transform 1 0 4312 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_28
timestamp 1663361622
transform 1 0 4468 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_29
timestamp 1663361622
transform 1 0 4624 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_30
timestamp 1663361622
transform 1 0 4780 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_31
timestamp 1663361622
transform 1 0 4936 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_32
timestamp 1663361622
transform 1 0 5092 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_33
timestamp 1663361622
transform 1 0 5248 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_34
timestamp 1663361622
transform 1 0 5404 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_35
timestamp 1663361622
transform 1 0 5560 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_36
timestamp 1663361622
transform 1 0 5716 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_37
timestamp 1663361622
transform 1 0 5872 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_38
timestamp 1663361622
transform 1 0 6028 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_39
timestamp 1663361622
transform 1 0 6184 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_40
timestamp 1663361622
transform 1 0 6340 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_41
timestamp 1663361622
transform 1 0 6496 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_42
timestamp 1663361622
transform 1 0 6652 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_43
timestamp 1663361622
transform 1 0 6808 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_44
timestamp 1663361622
transform 1 0 6964 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_45
timestamp 1663361622
transform 1 0 7120 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_46
timestamp 1663361622
transform 1 0 7276 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_47
timestamp 1663361622
transform 1 0 7432 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_48
timestamp 1663361622
transform 1 0 7588 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808336  sky130_fd_pr__dfl1sd__example_55959141808336_0
timestamp 1663361622
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808336  sky130_fd_pr__dfl1sd__example_55959141808336_1
timestamp 1663361622
transform 1 0 7744 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 11874496
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 11848162
<< end >>
