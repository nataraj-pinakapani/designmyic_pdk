magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 57 23 60 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 53 0 56 27 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 52 21 55 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 48 0 51 21 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 52 23 61 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 41 1 44 4 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 52 20 52 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 41 1 44 4 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 56 22 57 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 60 23 61 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 37 0 40 1 8 VSSA
port 3 nsew ground bidirectional
rlabel  s 48 0 57 27 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 56 0 57 27 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 52 0 53 22 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 37 0 40 1 8 VSSA
port 3 nsew ground bidirectional
rlabel  s 48 0 48 24 6 VSSA
port 3 nsew ground bidirectional
rlabel  s 0 19 1 22 4 VDDA
port 4 nsew power bidirectional
rlabel  s 0 19 1 22 4 VDDA
port 4 nsew power bidirectional
rlabel  s 15 0 18 1 8 VDDA
port 4 nsew power bidirectional
rlabel  s 15 0 18 1 8 VDDA
port 4 nsew power bidirectional
rlabel  s 0 36 1 39 4 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 36 1 39 4 VSWITCH
port 5 nsew power bidirectional
rlabel  s 32 0 35 1 8 VSWITCH
port 5 nsew power bidirectional
rlabel  s 32 0 35 1 8 VSWITCH
port 5 nsew power bidirectional
rlabel  s 0 68 1 72 4 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 68 1 73 4 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 64 0 68 1 8 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 64 0 69 1 8 VDDIO_Q
port 6 nsew power bidirectional
rlabel  s 0 6 2 11 6 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 6 2 11 6 VCCHIB
port 7 nsew power bidirectional
rlabel  s 2 0 7 1 8 VCCHIB
port 7 nsew power bidirectional
rlabel  s 2 0 7 1 8 VCCHIB
port 7 nsew power bidirectional
rlabel  s 0 74 3 99 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 24 2 28 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 24 2 28 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 74 3 99 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 20 0 24 1 8 VDDIO
port 8 nsew power bidirectional
rlabel  s 70 0 95 2 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 70 0 95 2 6 VDDIO
port 8 nsew power bidirectional
rlabel  s 20 0 24 1 8 VDDIO
port 8 nsew power bidirectional
rlabel  s 0 13 4 17 6 VCCD
port 9 nsew power bidirectional
rlabel  s 0 13 4 18 6 VCCD
port 9 nsew power bidirectional
rlabel  s 9 0 13 1 8 VCCD
port 9 nsew power bidirectional
rlabel  s 9 0 14 1 8 VCCD
port 9 nsew power bidirectional
rlabel  s 0 30 2 34 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 30 2 34 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 180 1 204 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 26 0 30 1 8 VSSIO
port 10 nsew ground bidirectional
rlabel  s 26 0 30 1 8 VSSIO
port 10 nsew ground bidirectional
rlabel  s 176 0 200 1 8 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 46 1 50 4 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 46 1 50 4 VSSD
port 11 nsew ground bidirectional
rlabel  s 42 0 46 1 8 VSSD
port 11 nsew ground bidirectional
rlabel  s 42 0 46 1 8 VSSD
port 11 nsew ground bidirectional
rlabel  s 0 62 2 67 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 62 2 67 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 58 0 63 1 8 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 58 0 63 1 8 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string LEFclass ENDCAP TOPRIGHT
string FIXED_BBOX 0 0 200 204
string LEFview TRUE
<< end >>
