magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal default
rlabel  s 79 53 80 56 6 AMUXBUS_A
port 1 nsew signal default
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal default
rlabel  s 79 48 80 51 6 AMUXBUS_B
port 2 nsew signal default
rlabel  s 32 128 53 149 6 PAD
port 3 nsew signal default
rlabel  s 79 13 80 14 6 VCCD
port 4 nsew power bidirectional
rlabel  s 79 9 80 9 6 VCCD
port 4 nsew power bidirectional
rlabel  s 0 13 1 14 4 VCCD
port 4 nsew power bidirectional
rlabel  s 0 9 80 13 6 VCCD
port 4 nsew power bidirectional
rlabel  s 0 9 1 9 4 VCCD
port 4 nsew power bidirectional
rlabel  s 0 9 80 13 6 VCCD
port 4 nsew power bidirectional
rlabel  s 79 7 80 7 6 VCCHIB
port 5 nsew power bidirectional
rlabel  s 79 2 80 2 6 VCCHIB
port 5 nsew power bidirectional
rlabel  s 0 7 1 7 4 VCCHIB
port 5 nsew power bidirectional
rlabel  s 0 2 80 7 6 VCCHIB
port 5 nsew power bidirectional
rlabel  s 0 2 1 2 4 VCCHIB
port 5 nsew power bidirectional
rlabel  s 0 2 80 7 6 VCCHIB
port 5 nsew power bidirectional
rlabel  s 0 18 1 18 4 VDDA
port 6 nsew power bidirectional
rlabel  s 0 15 79 18 6 VDDA
port 6 nsew power bidirectional
rlabel  s 0 15 1 15 4 VDDA
port 6 nsew power bidirectional
rlabel  s 79 15 80 18 6 VDDA
port 6 nsew power bidirectional
rlabel  s 0 15 80 18 6 VDDA
port 6 nsew power bidirectional
rlabel  s 79 24 80 24 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 79 20 80 20 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 24 1 24 4 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 20 80 24 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 20 1 20 4 VDDIO
port 7 nsew power bidirectional
rlabel  s 79 95 80 95 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 79 70 80 70 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 95 1 95 4 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 70 80 95 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 70 1 70 4 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 20 80 24 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 0 70 80 95 6 VDDIO
port 7 nsew power bidirectional
rlabel  s 79 68 80 69 6 VDDIO_Q
port 8 nsew power bidirectional
rlabel  s 79 64 80 64 6 VDDIO_Q
port 8 nsew power bidirectional
rlabel  s 0 68 1 69 4 VDDIO_Q
port 8 nsew power bidirectional
rlabel  s 0 64 80 68 6 VDDIO_Q
port 8 nsew power bidirectional
rlabel  s 0 64 1 64 4 VDDIO_Q
port 8 nsew power bidirectional
rlabel  s 0 64 80 68 6 VDDIO_Q
port 8 nsew power bidirectional
rlabel  s 79 40 80 40 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 79 37 80 37 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 40 1 40 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 37 80 40 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 37 1 37 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 48 1 48 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 52 80 53 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 56 1 57 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 79 48 80 48 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 79 56 80 57 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 37 80 40 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 48 80 57 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 79 46 80 46 6 VSSD
port 10 nsew ground bidirectional
rlabel  s 79 42 80 42 6 VSSD
port 10 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSD
port 10 nsew ground bidirectional
rlabel  s 0 42 80 46 6 VSSD
port 10 nsew ground bidirectional
rlabel  s 0 42 1 42 4 VSSD
port 10 nsew ground bidirectional
rlabel  s 0 42 80 46 6 VSSD
port 10 nsew ground bidirectional
rlabel  s 79 200 80 200 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 79 176 80 176 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 200 1 200 4 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 176 80 200 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 176 1 176 4 VSSIO
port 11 nsew ground bidirectional
rlabel  s 79 30 80 30 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 79 26 80 26 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 30 1 30 4 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 26 80 30 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 26 1 26 4 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 176 80 200 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 0 26 80 30 6 VSSIO
port 11 nsew ground bidirectional
rlabel  s 79 62 80 63 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 79 58 80 58 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 62 1 63 4 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 58 80 62 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 58 1 58 4 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 0 58 80 63 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel  s 79 35 80 35 6 VSWITCH
port 13 nsew power bidirectional
rlabel  s 79 32 80 32 6 VSWITCH
port 13 nsew power bidirectional
rlabel  s 0 35 1 35 4 VSWITCH
port 13 nsew power bidirectional
rlabel  s 0 32 80 35 6 VSWITCH
port 13 nsew power bidirectional
rlabel  s 0 32 1 32 4 VSWITCH
port 13 nsew power bidirectional
rlabel  s 0 32 80 35 6 VSWITCH
port 13 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 80 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
