magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel 
 s 26 0 37 20 6 DRN_LVC1
port 3 nsew power bidirectional
rlabel 
 s 38 0 49 23 6 DRN_LVC2
port 4 nsew power bidirectional
rlabel � s 1 0 20 1 8 SRC_BDY_LVC1
port 5 nsew ground bidirectional
rlabel � s 55 0 75 4 6 SRC_BDY_LVC2
port 6 nsew ground bidirectional
rlabel � s 34 0 44 0 8 BDY2_B2B
port 7 nsew ground bidirectional
rlabel  s 10 100 65 167 6 VDDIO_PAD
port 8 nsew power bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 54 75 55 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 46 75 46 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 9 nsew ground bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 10 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 10 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 10 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 10 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 11 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 11 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 11 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 11 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 13 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 13 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 13 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 13 nsew power bidirectional
rlabel 
 s 51 0 75 18 6 VDDIO
port 14 nsew power bidirectional
rlabel 
 s 1 0 25 18 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 14 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 15 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 15 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 15 nsew power bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 15 nsew power bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 16 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 16 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 16 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 16 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 16 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 16 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 17 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 17 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 17 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 17 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 18 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 18 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 18 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 18 nsew ground bidirectional
<< properties >>
string LEFclass PAD POWER
string FIXED_BBOX 0 0 75 198
string LEFview TRUE
<< end >>
