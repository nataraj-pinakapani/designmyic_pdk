magic
tech minimum
timestamp 1644097874
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -6 -3 7 18
string LEFview TRUE
<< end >>
