magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 53 75 56 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 48 75 51 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 37 139 38 146 6 G_PAD
port 3 nsew signal bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 175 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 175 74 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 152 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 152 74 152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 129 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 129 74 129 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 106 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 106 74 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 83 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 83 74 83 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 60 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 60 74 60 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 31 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 31 74 31 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 60 74 60 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 175 74 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 31 74 31 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 152 74 152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 129 74 129 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 106 74 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 83 74 83 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 60 74 60 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 175 74 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 31 74 31 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 152 74 152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 129 74 129 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 106 74 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 83 74 83 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 60 74 60 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 174 74 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 31 74 31 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 152 74 152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 128 74 129 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 105 74 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 82 74 83 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 59 74 60 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 31 74 31 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 151 74 152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 31 74 31 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 30 74 31 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 183 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 90 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 183 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 159 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 136 74 136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 113 74 113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 90 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 67 74 67 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 44 74 44 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 61 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 136 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 113 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 67 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 44 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 174 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 128 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 105 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 82 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 59 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 173 74 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 151 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 127 74 128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 104 74 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 81 74 82 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 58 74 59 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 150 74 151 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 30 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 29 74 30 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 91 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 137 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 91 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 68 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 45 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 184 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 160 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 137 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 114 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 68 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 60 45 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 173 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 127 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 104 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 81 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 58 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 172 74 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 150 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 126 74 127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 103 74 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 80 74 81 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 57 74 58 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 149 74 150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 29 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 185 74 185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 28 74 29 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 92 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 92 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 69 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 161 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 138 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 115 74 115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 69 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 46 74 46 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 59 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 115 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 46 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 172 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 126 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 103 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 80 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 57 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 171 74 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 149 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 125 74 126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 102 74 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 79 74 80 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 56 74 57 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 171 74 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 148 74 149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 125 74 125 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 102 74 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 79 74 79 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 171 74 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 28 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 125 74 125 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 102 74 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 79 74 79 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 171 74 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 27 74 28 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 125 74 125 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 102 74 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 79 74 79 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 171 74 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 125 74 125 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 102 74 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 79 74 79 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 93 74 93 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 162 74 162 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 139 74 139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 116 74 116 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 70 74 70 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 58 47 74 47 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 27 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 26 74 27 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 57 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 56 26 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 0 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 9 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 50 9 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 10 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 10 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 49 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 11 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 48 11 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 47 12 74 12 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 38 12 74 26 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 116 74 125 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 93 74 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 76 74 79 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 76 74 76 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 73 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 70 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 76 74 76 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 73 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 75 74 76 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 73 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 73 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 73 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 25 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 73 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 73 74 73 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 73 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 75 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 75 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 24 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 19 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 19 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 19 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 19 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 19 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 19 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 74 74 74 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 56 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 56 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 148 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 147 74 148 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 55 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 18 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 147 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 162 74 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 139 74 147 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 17 47 74 55 6 DRN_HVC
port 4 nsew power bidirectional
rlabel � s 16 185 74 190 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 169 59 169 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 110 59 169 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 110 59 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 110 59 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 169 59 169 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 110 59 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 169 59 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 110 59 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 170 59 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 110 59 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 170 59 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 110 59 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 53 170 59 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 109 59 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 170 59 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 109 59 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 170 59 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 109 59 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 170 59 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 109 59 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 170 59 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 109 59 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 171 59 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 109 59 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 171 59 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 52 109 59 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 171 59 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 108 59 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 171 59 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 108 59 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 171 59 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 108 59 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 171 59 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 108 59 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 172 59 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 108 59 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 172 59 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 108 59 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 172 59 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 51 108 59 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 172 59 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 107 59 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 172 59 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 107 59 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 172 59 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 107 58 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 172 59 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 107 58 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 173 59 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 175 61 190 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 175 61 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 175 61 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 174 61 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 174 60 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 174 60 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 174 60 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 174 60 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 174 60 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 173 60 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 173 60 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 173 59 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 173 59 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 173 59 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 107 58 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 50 107 58 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 49 106 58 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 49 106 58 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 49 106 57 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 49 106 57 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 49 106 57 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 49 106 57 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 49 106 57 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 48 105 57 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 48 105 57 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 48 105 56 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 48 105 56 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 48 105 56 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 48 105 56 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 48 105 56 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 47 104 56 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 47 104 56 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 47 104 55 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 47 104 55 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 47 104 55 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 47 104 55 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 46 103 55 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 46 103 55 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 46 103 54 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 46 103 54 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 46 103 54 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 46 103 54 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 46 103 54 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 102 54 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 102 54 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 102 53 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 102 53 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 102 53 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 102 53 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 102 53 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 101 53 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 101 53 101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 101 52 101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 101 52 101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 101 52 101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 101 52 101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 101 52 101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 52 101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 52 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 51 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 51 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 51 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 51 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 51 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 45 100 51 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 43 170 49 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 43 111 49 170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 43 111 49 111 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 43 110 49 111 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 43 171 49 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 43 110 49 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 43 171 49 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 110 49 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 171 49 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 110 49 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 171 49 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 110 49 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 171 49 171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 110 49 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 171 49 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 110 49 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 172 49 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 109 49 110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 172 49 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 109 49 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 42 172 49 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 109 49 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 172 49 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 109 49 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 172 49 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 109 49 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 172 49 172 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 109 49 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 172 49 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 108 49 109 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 173 49 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 108 49 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 173 49 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 41 108 49 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 173 49 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 108 49 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 173 49 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 108 49 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 173 49 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 108 48 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 173 49 173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 108 48 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 173 49 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 107 48 108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 174 49 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 107 48 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 174 49 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 40 107 48 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 174 49 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 107 48 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 174 49 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 107 48 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 174 49 174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 107 47 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 174 49 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 107 47 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 175 49 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 106 47 107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 175 49 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 106 47 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 39 175 49 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 106 47 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 175 49 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 106 47 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 175 49 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 106 47 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 175 49 175 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 106 46 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 175 49 190 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 106 46 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 105 46 106 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 105 46 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 105 46 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 105 46 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 105 46 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 105 45 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 105 45 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 104 45 105 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 104 45 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 104 45 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 104 45 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 104 44 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 104 44 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 103 44 104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 103 44 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 103 44 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 103 44 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 103 44 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 103 43 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 103 43 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 102 43 103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 102 43 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 102 43 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 100 43 102 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 100 43 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 100 43 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 100 43 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 100 43 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 100 43 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 98 51 100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 98 51 98 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 98 51 98 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 98 51 98 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 98 51 98 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 98 50 98 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 98 50 98 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 97 50 98 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 97 50 97 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 97 50 97 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 97 50 97 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 97 49 97 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 97 49 97 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 96 49 97 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 96 49 96 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 96 49 96 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 38 0 49 96 6 DRN_HVC
port 4 nsew power bidirectional
rlabel 
 s 1 46 24 47 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 37 24 46 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 37 24 37 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 37 24 37 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 47 24 47 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 37 24 37 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 47 24 47 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 37 24 37 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 1 47 24 47 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 101 14 173 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 101 14 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 101 14 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 101 14 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 101 14 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 101 14 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 101 14 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 100 14 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 100 14 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 100 15 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 100 15 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 100 15 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 100 15 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 100 15 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 99 15 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 99 16 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 99 16 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 99 16 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 99 16 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 99 16 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 98 16 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 98 16 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 98 17 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 98 17 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 98 17 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 98 17 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 98 17 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 97 17 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 97 17 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 97 18 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 97 18 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 97 18 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 97 18 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 97 18 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 96 18 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 96 19 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 96 19 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 96 19 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 96 19 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 96 19 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 95 19 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 95 19 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 95 20 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 95 20 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 95 20 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 95 20 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 95 20 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 94 20 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 94 20 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 94 21 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 94 21 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 94 21 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 94 21 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 94 21 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 93 21 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 93 22 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 93 22 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 93 22 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 93 22 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 93 22 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 92 22 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 92 22 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 92 23 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 92 23 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 92 23 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 92 23 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 92 23 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 91 23 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 91 23 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 91 24 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 91 24 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 91 24 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 91 24 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 91 24 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 47 24 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 0 0 24 37 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 62 101 74 173 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 62 101 74 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 61 101 74 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 61 101 74 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 61 101 74 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 61 101 74 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 61 101 74 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 61 100 74 101 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 61 100 74 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 60 100 74 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 60 100 74 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 60 100 74 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 60 100 74 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 60 99 74 100 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 60 99 74 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 60 99 74 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 59 99 74 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 59 99 74 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 59 99 74 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 59 99 74 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 59 98 74 99 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 59 98 74 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 58 98 74 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 58 98 74 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 58 98 74 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 58 98 74 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 58 98 74 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 58 97 74 98 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 58 97 74 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 57 97 74 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 57 97 74 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 57 97 74 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 57 97 74 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 57 96 74 97 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 57 96 74 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 57 96 74 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 56 96 74 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 56 96 74 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 56 96 74 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 56 96 74 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 56 95 74 96 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 56 95 74 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 55 95 74 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 55 95 74 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 55 95 74 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 55 95 74 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 55 95 74 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 55 94 74 95 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 55 94 74 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 54 94 74 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 54 94 74 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 54 94 74 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 54 94 74 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 54 93 74 94 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 54 93 74 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 54 93 74 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 53 93 74 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 53 93 74 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 53 93 74 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 53 93 74 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 53 92 74 93 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 53 92 74 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 52 92 74 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 52 92 74 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 52 92 74 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 52 92 74 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 52 92 74 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 52 91 74 92 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 52 91 74 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 51 91 74 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 51 91 74 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 51 91 74 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 51 91 74 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 51 90 74 91 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 51 90 74 90 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 51 90 74 90 6 G_CORE
port 5 nsew ground bidirectional
rlabel 
 s 50 0 74 90 6 G_CORE
port 5 nsew ground bidirectional
rlabel � s 26 0 28 1 8 OGC_HVC
port 6 nsew power bidirectional
rlabel � s 55 38 57 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 55 36 57 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 55 38 57 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 55 38 57 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 38 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 54 39 57 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 39 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 57 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 56 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 56 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 56 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 56 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 53 40 56 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 47 14 47 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 14 47 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 14 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 14 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 14 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 14 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 14 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 14 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 15 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 15 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 15 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 15 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 45 15 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 45 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 15 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 16 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 16 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 16 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 16 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 16 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 44 16 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 44 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 16 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 17 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 17 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 17 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 17 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 43 17 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 17 43 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 17 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 54 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 54 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 54 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 54 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 54 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 42 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 55 42 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 55 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 55 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 55 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 55 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 55 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 55 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 41 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 56 41 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 56 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 56 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 20 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 20 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 20 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 20 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 20 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 40 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 40 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 19 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 18 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 18 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 18 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 18 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 18 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 39 18 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 39 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 18 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 17 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 17 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 17 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 17 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 17 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 38 17 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 38 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 17 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 47 14 47 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 47 14 47 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 191 67 195 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 191 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 15 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 190 14 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 14 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 185 15 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 185 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 15 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 16 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 184 16 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 184 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 16 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 17 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 183 17 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 183 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 17 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 182 18 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 181 18 182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 173 58 181 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 173 18 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 173 18 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 173 17 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 173 17 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 17 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 172 16 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 16 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 171 15 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 15 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 170 14 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 169 14 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 169 14 169 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 169 14 169 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 169 14 169 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 14 169 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 14 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 14 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 14 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 14 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 14 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 14 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 15 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 162 15 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 15 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 16 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 161 16 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 16 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 17 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 160 17 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 17 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 18 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 159 18 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 158 18 159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 150 57 158 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 150 18 150 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 150 18 150 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 150 17 150 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 150 17 150 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 150 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 17 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 149 16 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 149 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 16 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 148 15 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 15 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 147 14 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 146 14 147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 146 14 146 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 146 14 146 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 146 14 146 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 146 14 146 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 14 146 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 14 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 14 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 14 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 14 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 14 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 14 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 15 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 15 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 139 15 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 15 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 16 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 16 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 16 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 138 16 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 16 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 17 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 17 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 137 17 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 17 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 18 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 18 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 136 18 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 135 18 136 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 127 57 135 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 127 18 127 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 127 18 127 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 127 18 127 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 127 17 127 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 127 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 126 17 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 125 16 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 124 15 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 123 14 124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 123 14 123 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 123 14 123 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 123 14 123 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 123 14 123 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 123 14 123 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 123 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 14 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 116 15 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 15 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 16 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 115 16 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 115 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 16 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 17 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 114 17 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 17 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 113 18 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 112 18 113 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 104 57 112 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 104 18 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 104 18 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 104 17 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 104 17 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 17 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 103 16 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 16 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 15 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 102 15 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 15 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 14 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 101 14 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 100 14 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 100 14 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 100 14 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 100 14 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 14 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 14 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 14 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 14 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 14 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 14 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 14 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 93 15 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 15 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 92 16 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 16 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 91 17 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 17 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 90 18 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 89 18 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 81 57 89 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 81 18 81 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 81 18 81 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 81 17 81 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 81 17 81 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 81 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 17 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 80 16 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 80 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 16 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 15 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 79 15 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 79 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 15 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 14 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 78 14 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 77 14 78 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 77 14 77 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 77 14 77 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 77 14 77 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 14 77 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 14 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 14 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 14 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 14 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 14 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 14 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 70 15 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 70 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 15 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 69 16 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 69 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 16 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 68 17 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 68 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 17 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 67 18 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 66 18 67 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 58 57 66 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 58 18 58 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 58 18 58 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 58 17 58 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 58 17 58 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 58 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 17 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 57 16 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 57 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 16 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 56 15 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 56 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 15 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 55 14 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 54 14 55 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 54 14 54 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 54 14 54 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 54 14 54 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 54 14 54 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 47 14 54 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 37 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 16 37 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 16 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 16 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 16 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 16 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 16 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 16 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 15 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 15 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 15 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 15 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 36 15 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 15 36 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 15 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 15 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 15 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 15 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 15 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 29 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 16 29 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 16 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 16 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 16 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 16 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 16 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 16 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 28 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 28 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 17 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 18 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 18 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 18 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 18 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 18 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 27 18 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 27 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 18 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 19 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 19 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 19 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 26 19 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 37 26 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 28 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 27 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 27 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 12 27 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 12 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 27 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 26 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 26 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 11 26 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 11 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 26 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 25 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 25 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 10 25 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 10 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 25 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 24 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 9 24 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 3 24 9 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 3 24 3 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 2 24 3 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 2 24 2 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 2 24 2 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 2 24 2 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 2 24 2 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 2 24 2 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 1 2 24 2 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel � s 0 0 24 2 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 96 37 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 93 37 96 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 93 37 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 93 37 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 97 37 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 93 37 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 97 37 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 32 93 37 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 97 37 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 92 37 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 97 37 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 97 37 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 97 37 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 97 37 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 98 37 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 31 98 37 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 30 98 37 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 30 98 37 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 30 98 37 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 30 98 37 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 30 98 37 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 30 99 37 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 30 99 37 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 29 99 37 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 29 99 37 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 29 99 37 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 29 99 37 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 29 100 37 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 29 100 37 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 100 37 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 100 37 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 100 37 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 100 36 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 100 36 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 100 36 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 101 36 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 28 101 36 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 27 101 36 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 27 101 36 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 27 101 35 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 27 101 35 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 27 102 35 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 27 102 35 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 102 35 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 102 35 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 102 34 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 102 34 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 175 37 195 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 175 37 175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 175 37 175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 175 36 175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 175 36 175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 175 36 175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 175 36 175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 174 36 175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 174 36 174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 174 36 174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 174 35 174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 174 35 174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 174 35 174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 173 35 174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 173 35 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 173 35 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 173 34 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 173 34 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 173 34 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 173 34 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 172 34 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 172 34 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 172 34 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 172 33 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 172 33 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 172 33 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 172 33 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 171 33 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 171 33 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 171 33 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 171 32 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 171 32 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 171 32 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 170 32 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 105 32 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 105 32 105 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 105 32 105 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 104 32 105 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 104 32 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 104 32 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 104 33 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 104 33 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 104 33 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 104 33 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 103 33 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 103 33 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 103 34 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 103 34 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 103 34 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 103 34 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 103 34 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 102 34 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 90 37 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 0 37 90 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 91 37 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 26 91 37 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 25 91 37 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 25 91 37 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 25 91 37 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 25 91 37 91 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 25 91 37 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 25 92 37 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 25 92 37 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 92 37 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 92 37 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 92 37 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 92 37 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 92 30 92 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 92 30 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 94 30 94 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 93 30 94 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 93 30 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 93 30 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 93 30 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 93 30 93 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 24 94 30 94 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 23 94 30 94 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 23 94 30 95 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 23 95 30 95 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 23 95 30 95 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 23 95 30 95 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 23 95 30 95 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 23 95 30 95 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 22 95 30 95 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 22 95 30 96 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 22 96 30 96 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 22 96 30 96 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 22 96 30 96 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 22 96 30 96 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 21 96 30 96 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 21 96 30 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 21 97 30 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 21 97 29 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 21 97 29 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 21 97 29 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 21 97 29 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 20 97 29 97 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 20 97 29 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 20 98 28 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 20 98 28 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 20 98 28 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 20 98 28 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 20 98 28 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 19 98 28 98 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 19 98 28 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 19 99 27 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 19 99 27 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 19 99 27 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 19 99 27 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 18 99 27 99 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 18 99 27 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 18 100 27 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 18 100 26 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 18 100 26 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 18 100 26 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 18 100 26 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 17 100 26 100 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 17 100 26 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 17 101 25 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 17 101 25 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 17 101 25 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 17 101 25 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 17 101 25 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 101 25 101 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 101 25 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 102 24 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 102 24 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 102 24 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 102 24 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 171 24 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 171 24 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 171 23 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 171 23 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 171 23 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 171 23 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 170 23 171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 170 23 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 170 23 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 170 22 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 170 22 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 170 22 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 170 22 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 169 22 170 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 169 22 169 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 169 22 169 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 105 22 169 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 105 22 105 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 104 22 105 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 104 22 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 104 22 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 104 22 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 104 22 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 104 22 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 104 22 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 103 23 104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 103 23 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 103 23 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 103 23 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 103 23 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 103 23 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 103 24 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 102 24 103 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 16 102 24 102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 15 171 24 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 15 172 24 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 15 172 24 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 15 172 24 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 15 172 24 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 15 172 25 172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 14 172 25 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 14 173 25 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 14 173 25 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 14 173 25 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 14 173 25 173 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel 
 s 14 173 25 195 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel  s 0 9 1 14 4 VCCD
port 8 nsew power bidirectional
rlabel  s 74 9 75 14 6 VCCD
port 8 nsew power bidirectional
rlabel  s 0 9 1 13 4 VCCD
port 8 nsew power bidirectional
rlabel  s 74 9 75 13 6 VCCD
port 8 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 9 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 9 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 9 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 9 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 10 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 10 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 10 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 10 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 11 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 74 64 75 69 6 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 0 64 1 68 4 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 74 64 75 68 6 VDDIO_Q
port 12 nsew power bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 13 nsew ground bidirectional
rlabel  s 0 48 1 48 4 VSSA
port 13 nsew ground bidirectional
rlabel  s 0 52 1 53 4 VSSA
port 13 nsew ground bidirectional
rlabel  s 0 56 1 57 4 VSSA
port 13 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 13 nsew ground bidirectional
rlabel  s 74 48 75 48 6 VSSA
port 13 nsew ground bidirectional
rlabel  s 74 52 75 53 6 VSSA
port 13 nsew ground bidirectional
rlabel  s 74 56 75 57 6 VSSA
port 13 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 13 nsew ground bidirectional
rlabel  s 0 48 1 57 4 VSSA
port 13 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 13 nsew ground bidirectional
rlabel  s 74 48 75 57 6 VSSA
port 13 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 14 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 14 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 14 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 14 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 15 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 15 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 15 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 15 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 15 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 15 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 15 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 15 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 16 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 16 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 17 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 17 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 17 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 17 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
