/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__esd_rf_diode_pw2nd_11v0_100__parasitic__diode_pw2dn.model.spice