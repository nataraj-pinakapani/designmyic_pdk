/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/fixed_devices/sky130_fd_pr__npn_05v5_W1p00L1p00_fail.cdl