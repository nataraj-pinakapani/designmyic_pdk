magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 79 53 80 56 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 79 48 80 51 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 62 0 63 2 6 ANALOG_EN
port 3 nsew signal input
rlabel 
 s 48 37 49 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 36 49 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 36 49 36 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 36 49 36 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 36 49 36 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 37 49 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 36 49 36 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 37 48 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 37 48 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 36 49 36 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 48 37 48 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 48 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 48 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 48 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 47 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 46 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 46 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 46 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 37 46 37 6 ANALOG_POL
port 4 nsew signal input
rlabel 
 s 46 0 46 37 6 ANALOG_POL
port 4 nsew signal input
rlabel � s 32 16 32 16 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 5 32 16 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 5 32 5 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 16 32 16 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 5 32 5 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 16 32 16 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 5 32 5 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 5 32 5 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 32 16 32 16 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 5 32 5 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 16 32 16 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 4 32 5 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 16 32 16 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 4 32 4 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 4 32 4 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 3 32 4 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 3 32 3 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 16 32 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 3 32 3 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 32 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 3 32 3 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 3 31 3 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 3 31 3 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 2 31 3 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 2 31 2 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 2 31 2 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 2 31 2 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 2 31 2 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 2 31 2 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 0 31 2 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 31 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 31 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 37 31 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 37 31 37 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 17 31 17 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 31 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 37 31 37 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 17 31 18 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 31 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 37 31 37 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 37 31 37 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 18 31 18 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 31 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 36 30 37 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 18 30 18 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 30 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 51 30 51 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 30 51 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 30 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 38 30 38 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 36 30 36 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 36 30 36 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 18 30 36 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 18 30 18 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 18 30 18 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 51 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 30 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 30 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 26 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 26 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 26 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 26 52 26 52 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 52 26 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 26 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 26 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 26 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 53 25 53 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 25 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 24 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 24 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 24 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 24 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 23 58 24 58 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 23 58 24 58 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 23 57 25 58 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 23 57 25 57 6 ANALOG_SEL
port 5 nsew signal input
rlabel � s 50 0 50 0 8 DM[0]
port 6 nsew signal input
rlabel � s 50 0 50 0 8 DM[0]
port 6 nsew signal input
rlabel � s 50 0 50 0 8 DM[0]
port 6 nsew signal input
rlabel � s 50 0 50 0 8 DM[0]
port 6 nsew signal input
rlabel � s 50 0 50 0 8 DM[0]
port 6 nsew signal input
rlabel � s 50 0 50 1 8 DM[0]
port 6 nsew signal input
rlabel � s 50 1 50 1 6 DM[0]
port 6 nsew signal input
rlabel � s 50 1 50 1 6 DM[0]
port 6 nsew signal input
rlabel � s 67 1 67 1 6 DM[1]
port 7 nsew signal input
rlabel � s 67 0 67 1 8 DM[1]
port 7 nsew signal input
rlabel � s 67 1 67 1 6 DM[1]
port 7 nsew signal input
rlabel � s 67 1 67 1 6 DM[1]
port 7 nsew signal input
rlabel � s 67 1 67 1 6 DM[1]
port 7 nsew signal input
rlabel � s 67 1 67 1 6 DM[1]
port 7 nsew signal input
rlabel � s 67 1 67 1 6 DM[1]
port 7 nsew signal input
rlabel � s 67 1 67 1 6 DM[1]
port 7 nsew signal input
rlabel � s 29 5 29 7 6 DM[2]
port 8 nsew signal input
rlabel � s 29 5 29 5 6 DM[2]
port 8 nsew signal input
rlabel � s 29 5 29 5 6 DM[2]
port 8 nsew signal input
rlabel � s 29 5 29 5 6 DM[2]
port 8 nsew signal input
rlabel � s 29 5 29 5 6 DM[2]
port 8 nsew signal input
rlabel � s 29 4 29 5 6 DM[2]
port 8 nsew signal input
rlabel � s 29 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 29 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 29 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 29 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 29 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 29 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 28 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 28 4 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 28 0 29 4 6 DM[2]
port 8 nsew signal input
rlabel � s 35 2 36 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 0 36 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 36 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 36 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 36 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 36 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 36 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 35 4 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 35 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 35 2 35 2 6 ENABLE_H
port 9 nsew signal input
rlabel � s 38 0 39 4 6 ENABLE_INP_H
port 10 nsew signal input
rlabel � s 15 32 16 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 20 16 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 20 16 20 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 16 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 20 16 20 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 16 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 16 20 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 16 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 16 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 15 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 15 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 15 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 37 15 37 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 15 37 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 15 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 32 15 32 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 37 15 37 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 37 15 37 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 37 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 15 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 19 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 18 15 19 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 15 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 18 14 18 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 14 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 18 14 18 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 14 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 18 14 18 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 14 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 18 14 18 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 18 14 18 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 7 14 18 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 7 14 7 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 14 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 6 14 7 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 14 38 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 38 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 14 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 14 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 6 14 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 13 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 6 13 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 13 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 6 13 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 13 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 6 13 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 13 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 5 13 6 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 13 39 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 5 13 5 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 39 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 5 13 5 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 5 13 5 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 5 13 5 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 0 13 5 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 13 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 13 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 12 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 12 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 12 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 12 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 12 40 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 40 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 12 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 12 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 11 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 11 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 11 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 11 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 11 41 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 41 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 11 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 11 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 10 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 10 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 10 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 10 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 10 42 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 42 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 10 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 10 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 9 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 9 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 9 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 9 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 9 43 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 43 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 9 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 77 8 77 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 77 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 54 8 54 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 8 54 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 8 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 44 9 44 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 77 8 77 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 54 8 54 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 77 8 77 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 77 9 77 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 54 8 54 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 54 8 54 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 54 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 54 8 54 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 54 8 54 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 77 9 78 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 75 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 74 8 75 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 8 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 56 8 56 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 74 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 57 8 74 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 57 8 57 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel � s 7 56 8 57 6 ENABLE_VDDA_H
port 11 nsew signal input
rlabel 
 s 79 0 79 176 6 ENABLE_VDDIO
port 12 nsew signal input
rlabel � s 18 37 18 37 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 18 36 18 37 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 18 35 18 36 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 18 37 18 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 18 35 18 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 18 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 18 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 18 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 18 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 18 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 18 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 18 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 18 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 18 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 35 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 31 17 31 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 12 17 31 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 12 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 7 17 7 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 3 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 34 17 35 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 38 17 38 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 31 17 31 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 2 17 3 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 34 17 34 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 17 31 17 31 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 38 17 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 2 17 2 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 34 17 34 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 31 17 32 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 17 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 2 17 2 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 32 17 32 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 34 17 34 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 34 17 34 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 32 17 34 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 32 17 32 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 32 17 32 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 17 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 2 17 2 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 2 17 2 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 0 17 2 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 17 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 17 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 39 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 16 39 16 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 15 40 16 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 15 40 16 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 16 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 58 15 58 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 58 15 58 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 58 15 58 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 49 15 58 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 49 15 49 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 16 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 49 15 49 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 58 15 58 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 15 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 49 15 49 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 48 15 49 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 58 15 58 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 58 15 58 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 15 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 41 14 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 41 14 41 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 41 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 40 14 40 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 42 14 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 14 42 14 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 14 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 14 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 14 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 14 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 42 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 42 13 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 13 43 13 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 13 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 13 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 13 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 13 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 14 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 43 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 12 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 12 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 43 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 12 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 44 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 12 48 12 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 44 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 48 12 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 44 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 47 12 48 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 44 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 47 12 47 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 44 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 47 12 47 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 47 12 47 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 44 12 47 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 44 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 11 44 12 44 6 ENABLE_VSWITCH_H
port 13 nsew signal input
rlabel � s 32 0 32 4 6 HLD_H_N
port 14 nsew signal input
rlabel � s 27 0 27 2 6 HLD_OVR
port 15 nsew signal input
rlabel � s 6 6 7 6 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 7 6 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 7 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 7 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 6 7 6 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 7 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 6 7 6 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 6 7 7 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 6 5 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 5 4 6 5 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 5 4 6 4 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 5 4 6 4 6 IB_MODE_SEL
port 16 nsew signal input
rlabel � s 5 0 6 4 6 IB_MODE_SEL
port 16 nsew signal input
rlabel 
 s 79 0 80 176 6 IN
port 17 nsew signal output
rlabel � s 46 6 46 7 6 INP_DIS
port 18 nsew signal input
rlabel � s 46 6 46 6 6 INP_DIS
port 18 nsew signal input
rlabel � s 46 6 46 6 6 INP_DIS
port 18 nsew signal input
rlabel � s 46 6 46 6 6 INP_DIS
port 18 nsew signal input
rlabel � s 46 6 46 6 6 INP_DIS
port 18 nsew signal input
rlabel � s 46 5 46 6 6 INP_DIS
port 18 nsew signal input
rlabel � s 46 5 46 5 6 INP_DIS
port 18 nsew signal input
rlabel � s 46 5 46 5 6 INP_DIS
port 18 nsew signal input
rlabel � s 45 5 46 5 6 INP_DIS
port 18 nsew signal input
rlabel � s 45 5 46 5 6 INP_DIS
port 18 nsew signal input
rlabel � s 45 5 46 5 6 INP_DIS
port 18 nsew signal input
rlabel � s 45 5 46 5 6 INP_DIS
port 18 nsew signal input
rlabel � s 45 5 46 5 6 INP_DIS
port 18 nsew signal input
rlabel � s 45 0 46 5 6 INP_DIS
port 18 nsew signal input
rlabel 
 s 3 181 5 181 6 IN_H
port 19 nsew signal output
rlabel 
 s 3 181 5 181 6 IN_H
port 19 nsew signal output
rlabel 
 s 3 181 5 181 6 IN_H
port 19 nsew signal output
rlabel 
 s 3 181 5 181 6 IN_H
port 19 nsew signal output
rlabel 
 s 3 180 5 181 6 IN_H
port 19 nsew signal output
rlabel 
 s 2 180 3 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 2 180 3 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 2 180 3 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 2 180 3 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 2 180 3 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 2 180 2 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 2 180 2 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 1 179 2 180 6 IN_H
port 19 nsew signal output
rlabel 
 s 1 179 2 179 6 IN_H
port 19 nsew signal output
rlabel 
 s 1 179 2 179 6 IN_H
port 19 nsew signal output
rlabel 
 s 1 179 2 179 6 IN_H
port 19 nsew signal output
rlabel 
 s 1 179 2 179 6 IN_H
port 19 nsew signal output
rlabel 
 s 1 179 1 179 6 IN_H
port 19 nsew signal output
rlabel 
 s 1 178 1 179 6 IN_H
port 19 nsew signal output
rlabel 
 s 0 178 1 178 4 IN_H
port 19 nsew signal output
rlabel 
 s 0 178 1 178 4 IN_H
port 19 nsew signal output
rlabel 
 s 0 0 1 178 4 IN_H
port 19 nsew signal output
rlabel � s 7 39 7 39 6 OE_N
port 20 nsew signal input
rlabel � s 7 10 7 39 6 OE_N
port 20 nsew signal input
rlabel � s 7 9 7 10 6 OE_N
port 20 nsew signal input
rlabel � s 7 39 7 39 6 OE_N
port 20 nsew signal input
rlabel � s 7 9 7 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 7 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 7 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 7 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 7 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 7 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 7 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 7 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 7 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 7 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 6 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 6 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 6 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 6 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 43 6 43 6 OE_N
port 20 nsew signal input
rlabel � s 6 43 6 43 6 OE_N
port 20 nsew signal input
rlabel � s 6 43 6 43 6 OE_N
port 20 nsew signal input
rlabel � s 6 40 6 43 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 6 40 6 OE_N
port 20 nsew signal input
rlabel � s 6 39 6 39 6 OE_N
port 20 nsew signal input
rlabel � s 6 43 6 43 6 OE_N
port 20 nsew signal input
rlabel � s 6 43 6 44 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 9 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 8 6 9 6 OE_N
port 20 nsew signal input
rlabel � s 6 8 6 8 6 OE_N
port 20 nsew signal input
rlabel � s 5 8 6 8 6 OE_N
port 20 nsew signal input
rlabel � s 5 8 6 8 6 OE_N
port 20 nsew signal input
rlabel � s 5 8 6 8 6 OE_N
port 20 nsew signal input
rlabel � s 5 5 6 8 6 OE_N
port 20 nsew signal input
rlabel � s 5 5 6 5 6 OE_N
port 20 nsew signal input
rlabel � s 5 5 6 5 6 OE_N
port 20 nsew signal input
rlabel � s 5 5 6 5 6 OE_N
port 20 nsew signal input
rlabel � s 5 5 6 5 6 OE_N
port 20 nsew signal input
rlabel � s 5 5 5 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 5 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 5 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 5 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 5 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 4 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 4 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 4 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 4 5 6 OE_N
port 20 nsew signal input
rlabel � s 4 5 4 5 6 OE_N
port 20 nsew signal input
rlabel � s 3 4 4 5 6 OE_N
port 20 nsew signal input
rlabel � s 3 4 4 4 6 OE_N
port 20 nsew signal input
rlabel � s 3 4 4 4 6 OE_N
port 20 nsew signal input
rlabel � s 3 0 4 4 6 OE_N
port 20 nsew signal input
rlabel � s 24 25 24 25 6 OUT
port 21 nsew signal input
rlabel � s 24 15 24 25 6 OUT
port 21 nsew signal input
rlabel � s 24 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 24 25 24 25 6 OUT
port 21 nsew signal input
rlabel � s 24 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 24 25 24 25 6 OUT
port 21 nsew signal input
rlabel � s 24 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 24 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 24 25 24 25 6 OUT
port 21 nsew signal input
rlabel � s 23 38 24 38 6 OUT
port 21 nsew signal input
rlabel � s 23 25 24 38 6 OUT
port 21 nsew signal input
rlabel � s 23 25 24 25 6 OUT
port 21 nsew signal input
rlabel � s 23 25 24 25 6 OUT
port 21 nsew signal input
rlabel � s 23 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 23 38 24 39 6 OUT
port 21 nsew signal input
rlabel � s 23 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 23 39 24 39 6 OUT
port 21 nsew signal input
rlabel � s 23 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 23 39 24 39 6 OUT
port 21 nsew signal input
rlabel � s 23 15 24 15 6 OUT
port 21 nsew signal input
rlabel � s 23 15 23 15 6 OUT
port 21 nsew signal input
rlabel � s 23 15 23 15 6 OUT
port 21 nsew signal input
rlabel � s 23 39 24 39 6 OUT
port 21 nsew signal input
rlabel � s 23 15 23 15 6 OUT
port 21 nsew signal input
rlabel � s 23 15 23 15 6 OUT
port 21 nsew signal input
rlabel � s 23 15 23 15 6 OUT
port 21 nsew signal input
rlabel � s 23 14 23 15 6 OUT
port 21 nsew signal input
rlabel � s 23 14 23 14 6 OUT
port 21 nsew signal input
rlabel � s 23 14 23 14 6 OUT
port 21 nsew signal input
rlabel � s 23 7 23 14 6 OUT
port 21 nsew signal input
rlabel � s 23 7 23 7 6 OUT
port 21 nsew signal input
rlabel � s 23 7 23 7 6 OUT
port 21 nsew signal input
rlabel � s 23 7 23 7 6 OUT
port 21 nsew signal input
rlabel � s 23 7 23 7 6 OUT
port 21 nsew signal input
rlabel � s 23 7 23 7 6 OUT
port 21 nsew signal input
rlabel � s 22 6 23 7 6 OUT
port 21 nsew signal input
rlabel � s 22 6 23 6 6 OUT
port 21 nsew signal input
rlabel � s 22 6 23 6 6 OUT
port 21 nsew signal input
rlabel � s 22 6 23 6 6 OUT
port 21 nsew signal input
rlabel � s 22 0 23 6 6 OUT
port 21 nsew signal input
rlabel  s 32 125 54 147 6 PAD
port 22 nsew signal bidirectional
rlabel � s 77 3 78 5 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 3 78 3 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 3 78 3 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 3 78 3 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 3 78 3 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 3 78 3 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 3 78 3 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 2 78 3 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 2 78 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 2 78 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 77 2 78 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 2 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 76 0 77 2 6 PAD_A_ESD_0_H
port 23 nsew signal bidirectional
rlabel � s 68 0 69 4 6 PAD_A_ESD_1_H
port 24 nsew signal bidirectional
rlabel 
 s 69 76 70 102 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 69 76 70 76 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 69 76 70 76 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 68 76 70 76 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 68 76 70 76 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 68 75 70 76 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 68 75 70 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 68 75 70 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 68 75 70 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 75 70 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 75 69 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 8 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 8 64 8 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 6 64 6 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 0 64 6 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 75 69 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 8 64 8 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 6 64 6 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 35 64 35 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 35 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 18 64 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 75 69 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 7 64 8 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 63 6 64 6 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 35 64 35 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 75 69 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 7 64 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 6 64 6 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 35 64 35 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 75 69 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 7 64 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 6 64 6 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 35 64 35 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 69 75 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 35 63 36 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 69 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 36 63 36 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 64 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 64 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 36 63 36 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 64 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 64 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 64 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 74 63 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 73 63 74 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 73 63 73 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 73 63 73 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 73 63 73 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 36 63 73 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 36 63 36 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 36 63 36 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 62 36 63 36 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 18 62 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 13 62 18 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 13 62 13 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 13 62 13 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 18 62 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 12 62 13 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 62 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 62 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 12 62 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 12 62 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 62 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 12 62 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 62 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 12 62 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 6 64 6 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 62 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 12 62 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 61 47 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 61 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 61 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 19 62 19 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 6 64 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 61 12 61 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 64 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 12 61 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 64 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 11 61 12 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 64 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 11 61 11 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 64 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 61 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 11 61 11 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 61 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 11 61 11 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 61 7 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 11 61 11 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 11 61 11 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 11 60 11 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 8 60 11 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 8 60 8 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 8 60 8 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel 
 s 60 7 61 8 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 10 121 13 121 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 10 105 13 105 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 10 121 13 121 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 10 105 13 105 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 10 121 13 121 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 10 105 13 105 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 121 13 121 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 105 13 105 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 121 13 121 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 105 13 105 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 120 13 121 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 105 13 106 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 120 13 120 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 106 13 106 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 120 13 120 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 106 13 106 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 120 13 120 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 106 13 106 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 9 120 13 120 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 106 13 106 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 120 13 120 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 106 13 106 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 120 13 120 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 106 13 106 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 119 13 120 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 106 13 107 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 119 13 119 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 107 13 107 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 119 13 119 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 8 119 13 119 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel  s 2 107 13 119 6 PAD_A_NOESD_H
port 25 nsew signal bidirectional
rlabel � s 78 1 78 1 6 SLOW
port 26 nsew signal input
rlabel � s 78 1 78 1 6 SLOW
port 26 nsew signal input
rlabel � s 78 1 78 1 6 SLOW
port 26 nsew signal input
rlabel � s 78 0 78 1 8 SLOW
port 26 nsew signal input
rlabel � s 78 1 78 1 6 SLOW
port 26 nsew signal input
rlabel � s 77 1 78 1 6 SLOW
port 26 nsew signal input
rlabel � s 77 1 78 1 6 SLOW
port 26 nsew signal input
rlabel � s 79 48 80 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 80 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 80 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 80 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 80 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 79 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 79 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 79 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 79 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 79 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 17 79 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 16 79 17 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 16 79 16 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 1 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 1 79 1 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 1 79 1 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 1 79 1 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 0 79 1 8 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 16 79 16 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 16 79 16 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 16 79 16 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 16 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 10 79 10 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 48 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 79 48 79 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 79 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 79 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 79 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 49 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 78 49 78 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 78 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 78 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 78 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 96 77 96 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 96 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 96 77 96 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 50 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 50 77 51 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 77 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 51 77 51 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 51 77 51 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 51 77 51 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 53 77 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 51 77 51 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 52 76 53 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 52 76 52 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 51 76 52 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 51 76 51 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 76 51 76 51 6 TIE_HI_ESD
port 27 nsew signal output
rlabel � s 80 0 80 96 6 TIE_LO_ESD
port 28 nsew signal output
rlabel � s 8 4 9 7 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 4 9 4 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 4 9 4 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 4 9 4 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 4 9 4 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 4 9 4 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 4 8 4 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 4 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 8 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 3 8 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 3 7 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 3 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 7 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 2 7 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 1 6 2 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 1 6 1 6 VTRIP_SEL
port 29 nsew signal input
rlabel � s 6 0 6 1 8 VTRIP_SEL
port 29 nsew signal input
rlabel  s 0 9 1 14 4 VCCD
port 30 nsew power bidirectional
rlabel  s 79 9 80 14 6 VCCD
port 30 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 31 nsew power bidirectional
rlabel  s 79 2 80 7 6 VCCHIB
port 31 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 32 nsew power bidirectional
rlabel  s 79 15 80 18 6 VDDA
port 32 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 33 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 33 nsew power bidirectional
rlabel  s 79 20 80 24 6 VDDIO
port 33 nsew power bidirectional
rlabel  s 79 70 80 95 6 VDDIO
port 33 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 34 nsew power bidirectional
rlabel  s 79 64 80 69 6 VDDIO_Q
port 34 nsew power bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 35 nsew ground bidirectional
rlabel  s 0 48 1 48 4 VSSA
port 35 nsew ground bidirectional
rlabel  s 0 52 1 53 4 VSSA
port 35 nsew ground bidirectional
rlabel  s 0 56 1 57 4 VSSA
port 35 nsew ground bidirectional
rlabel  s 79 37 80 40 6 VSSA
port 35 nsew ground bidirectional
rlabel  s 79 48 80 48 6 VSSA
port 35 nsew ground bidirectional
rlabel  s 79 52 80 53 6 VSSA
port 35 nsew ground bidirectional
rlabel  s 79 56 80 57 6 VSSA
port 35 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 36 nsew ground bidirectional
rlabel  s 79 42 80 46 6 VSSD
port 36 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 176 80 200 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 26 80 30 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 38 nsew ground bidirectional
rlabel  s 79 58 80 63 6 VSSIO_Q
port 38 nsew ground bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 39 nsew power bidirectional
rlabel  s 79 32 80 35 6 VSWITCH
port 39 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 80 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
