magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 5 4 5 9 6 BULK
port 1 nsew
rlabel  s 1 4 1 9 6 BULK
port 1 nsew
rlabel  s 0 5 6 8 6 DRAIN
port 2 nsew
rlabel  s 2 9 5 9 6 GATE
port 3 nsew
rlabel  s 2 3 5 3 6 GATE
port 3 nsew
rlabel  s 0 10 6 13 6 SOURCE
port 4 nsew
rlabel  s 0 0 6 3 6 SOURCE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 6 13
string LEFview TRUE
<< end >>
