magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 82 21 567 157
rect 29 -17 63 17
<< locali >>
rect 121 326 172 487
rect 293 326 344 487
rect 464 326 516 487
rect 21 292 627 326
rect 21 179 55 292
rect 89 213 532 258
rect 567 179 627 292
rect 21 145 627 179
rect 206 56 258 145
rect 378 56 429 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 360 86 527
rect 206 360 258 527
rect 378 360 430 527
rect 550 360 627 527
rect 113 17 172 111
rect 292 17 344 111
rect 463 17 523 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 89 213 532 258 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 378 56 429 145 6 Y
port 6 nsew signal output
rlabel locali s 206 56 258 145 6 Y
port 6 nsew signal output
rlabel locali s 21 145 627 179 6 Y
port 6 nsew signal output
rlabel locali s 567 179 627 292 6 Y
port 6 nsew signal output
rlabel locali s 21 179 55 292 6 Y
port 6 nsew signal output
rlabel locali s 21 292 627 326 6 Y
port 6 nsew signal output
rlabel locali s 464 326 516 487 6 Y
port 6 nsew signal output
rlabel locali s 293 326 344 487 6 Y
port 6 nsew signal output
rlabel locali s 121 326 172 487 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3365102
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3359296
<< end >>
