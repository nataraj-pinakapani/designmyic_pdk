magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 821 157 1195 203
rect 1 21 1195 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 538 47 568 131
rect 624 47 654 131
rect 711 47 741 131
rect 899 47 929 177
rect 995 47 1025 177
rect 1087 47 1117 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 530 425 560 497
rect 634 425 664 497
rect 747 413 777 497
rect 899 297 929 497
rect 995 297 1025 497
rect 1087 297 1117 497
<< ndiff >>
rect 847 161 899 177
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 47 538 131
rect 568 107 624 131
rect 568 73 579 107
rect 613 73 624 107
rect 568 47 624 73
rect 654 47 711 131
rect 741 106 793 131
rect 741 72 751 106
rect 785 72 793 106
rect 741 47 793 72
rect 847 127 855 161
rect 889 127 899 161
rect 847 93 899 127
rect 847 59 855 93
rect 889 59 899 93
rect 847 47 899 59
rect 929 47 995 177
rect 1025 127 1087 177
rect 1025 93 1043 127
rect 1077 93 1087 127
rect 1025 47 1087 93
rect 1117 133 1169 177
rect 1117 99 1127 133
rect 1161 99 1169 133
rect 1117 47 1169 99
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 425 530 497
rect 560 485 634 497
rect 560 451 578 485
rect 612 451 634 485
rect 560 425 634 451
rect 664 425 747 497
rect 465 369 515 425
rect 697 413 747 425
rect 777 477 899 497
rect 777 443 787 477
rect 821 443 855 477
rect 889 443 899 477
rect 777 413 899 443
rect 849 297 899 413
rect 929 471 995 497
rect 929 437 946 471
rect 980 437 995 471
rect 929 368 995 437
rect 929 334 946 368
rect 980 334 995 368
rect 929 297 995 334
rect 1025 485 1087 497
rect 1025 451 1043 485
rect 1077 451 1087 485
rect 1025 417 1087 451
rect 1025 383 1043 417
rect 1077 383 1087 417
rect 1025 297 1087 383
rect 1117 475 1169 497
rect 1117 441 1127 475
rect 1161 441 1169 475
rect 1117 384 1169 441
rect 1117 350 1127 384
rect 1161 350 1169 384
rect 1117 297 1169 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 579 73 613 107
rect 751 72 785 106
rect 855 127 889 161
rect 855 59 889 93
rect 1043 93 1077 127
rect 1127 99 1161 133
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 578 451 612 485
rect 787 443 821 477
rect 855 443 889 477
rect 946 437 980 471
rect 946 334 980 368
rect 1043 451 1077 485
rect 1043 383 1077 417
rect 1127 441 1161 475
rect 1127 350 1161 384
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 530 497 560 523
rect 634 497 664 523
rect 747 497 777 523
rect 899 497 929 523
rect 995 497 1025 523
rect 1087 497 1117 523
rect 79 348 109 363
rect 45 318 109 348
rect 45 280 75 318
rect 21 264 75 280
rect 163 274 193 363
rect 351 343 381 369
rect 21 230 31 264
rect 65 230 75 264
rect 21 214 75 230
rect 117 264 193 274
rect 117 230 133 264
rect 167 230 193 264
rect 317 313 381 343
rect 317 241 347 313
rect 117 220 193 230
rect 45 176 75 214
rect 45 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 293 225 381 241
rect 293 191 303 225
rect 337 191 381 225
rect 435 219 465 369
rect 530 338 560 425
rect 634 387 664 425
rect 603 377 669 387
rect 603 343 619 377
rect 653 343 669 377
rect 747 373 777 413
rect 530 337 561 338
rect 507 321 561 337
rect 603 333 669 343
rect 719 357 807 373
rect 507 287 517 321
rect 551 291 561 321
rect 719 323 763 357
rect 797 323 807 357
rect 719 307 807 323
rect 551 287 654 291
rect 507 261 654 287
rect 293 175 381 191
rect 351 131 381 175
rect 423 203 477 219
rect 423 169 433 203
rect 467 169 477 203
rect 423 153 477 169
rect 528 203 582 219
rect 528 169 538 203
rect 572 169 582 203
rect 528 153 582 169
rect 435 131 465 153
rect 538 131 568 153
rect 624 131 654 261
rect 719 181 749 307
rect 899 265 929 297
rect 995 265 1025 297
rect 1087 265 1117 297
rect 791 249 929 265
rect 791 215 801 249
rect 835 215 929 249
rect 791 199 929 215
rect 971 249 1025 265
rect 971 215 981 249
rect 1015 215 1025 249
rect 971 199 1025 215
rect 1067 249 1121 265
rect 1067 215 1077 249
rect 1111 215 1121 249
rect 1067 199 1121 215
rect 711 151 749 181
rect 899 177 929 199
rect 995 177 1025 199
rect 1087 177 1117 199
rect 711 131 741 151
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 538 21 568 47
rect 624 21 654 47
rect 711 21 741 47
rect 899 21 929 47
rect 995 21 1025 47
rect 1087 21 1117 47
<< polycont >>
rect 31 230 65 264
rect 133 230 167 264
rect 303 191 337 225
rect 619 343 653 377
rect 517 287 551 321
rect 763 323 797 357
rect 433 169 467 203
rect 538 169 572 203
rect 801 215 835 249
rect 981 215 1015 249
rect 1077 215 1111 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 247 493
rect 391 485 449 527
rect 237 443 247 477
rect 17 375 35 409
rect 203 409 247 443
rect 69 375 155 393
rect 17 359 155 375
rect 17 264 65 325
rect 17 230 31 264
rect 17 197 65 230
rect 121 323 155 359
rect 121 280 155 289
rect 237 391 247 409
rect 203 357 213 375
rect 203 337 247 357
rect 286 449 307 483
rect 341 449 357 483
rect 286 415 357 449
rect 286 381 307 415
rect 341 381 357 415
rect 121 264 167 280
rect 121 230 133 264
rect 121 214 167 230
rect 121 161 155 214
rect 34 127 155 161
rect 34 119 69 127
rect 34 85 35 119
rect 203 119 237 337
rect 286 333 357 381
rect 425 451 449 485
rect 562 451 578 485
rect 612 451 725 485
rect 391 417 449 451
rect 425 383 449 417
rect 391 367 449 383
rect 580 391 653 399
rect 580 357 585 391
rect 619 377 653 391
rect 601 343 619 357
rect 286 299 423 333
rect 287 225 353 265
rect 287 191 303 225
rect 337 191 353 225
rect 389 219 423 299
rect 489 325 552 337
rect 601 327 653 343
rect 489 323 567 325
rect 523 321 567 323
rect 489 287 517 289
rect 551 287 567 321
rect 489 271 567 287
rect 601 219 649 327
rect 691 265 725 451
rect 786 477 889 527
rect 786 443 787 477
rect 821 443 855 477
rect 786 427 889 443
rect 925 471 993 487
rect 925 437 946 471
rect 980 437 993 471
rect 925 373 993 437
rect 1027 485 1093 527
rect 1027 451 1043 485
rect 1077 451 1093 485
rect 1027 417 1093 451
rect 1027 383 1043 417
rect 1077 383 1093 417
rect 1127 475 1179 491
rect 1161 441 1179 475
rect 1127 384 1179 441
rect 763 368 993 373
rect 763 357 946 368
rect 797 334 946 357
rect 980 347 993 368
rect 1161 350 1179 384
rect 980 334 1093 347
rect 1127 334 1179 350
rect 797 323 1093 334
rect 763 307 1093 323
rect 869 301 1093 307
rect 691 249 835 265
rect 691 233 801 249
rect 389 203 467 219
rect 389 169 433 203
rect 389 157 467 169
rect 34 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 302 153 467 157
rect 538 203 649 219
rect 572 169 649 203
rect 538 153 649 169
rect 683 215 801 233
rect 683 199 835 215
rect 302 123 423 153
rect 302 119 341 123
rect 302 85 307 119
rect 683 107 717 199
rect 869 161 915 301
rect 1049 265 1093 301
rect 839 127 855 161
rect 889 127 915 161
rect 302 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 563 73 579 107
rect 613 73 717 107
rect 751 106 805 122
rect 375 17 441 55
rect 785 72 805 106
rect 751 17 805 72
rect 839 93 915 127
rect 839 59 855 93
rect 889 59 915 93
rect 949 249 1015 265
rect 949 215 981 249
rect 949 199 1015 215
rect 1049 249 1111 265
rect 1049 215 1077 249
rect 1049 199 1111 215
rect 949 69 995 199
rect 1145 149 1179 334
rect 1031 127 1088 143
rect 1031 93 1043 127
rect 1077 93 1088 127
rect 1031 17 1088 93
rect 1122 133 1179 149
rect 1122 99 1127 133
rect 1161 99 1179 133
rect 1122 69 1179 99
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 121 289 155 323
rect 213 375 237 391
rect 237 375 247 391
rect 213 357 247 375
rect 585 357 619 391
rect 489 321 523 323
rect 489 289 517 321
rect 517 289 523 321
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 573 391 631 397
rect 573 388 585 391
rect 247 360 585 388
rect 247 357 259 360
rect 201 351 259 357
rect 573 357 585 360
rect 619 357 631 391
rect 573 351 631 357
rect 109 323 167 329
rect 109 289 121 323
rect 155 320 167 323
rect 477 323 535 329
rect 477 320 489 323
rect 155 292 489 320
rect 155 289 167 292
rect 109 283 167 289
rect 477 289 489 292
rect 523 289 535 323
rect 477 283 535 289
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1133 357 1167 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1133 425 1167 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1133 85 1167 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 949 85 983 119 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 949 153 983 187 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlrtp_1
rlabel metal1 s 0 -48 1196 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 2786766
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 2776028
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 29.900 0.000 
<< end >>
