magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 53 1 56 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 53 75 56 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 48 1 51 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 48 75 51 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 9 1 14 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 9 75 14 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 9 1 13 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 9 75 13 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 4 nsew power bidirectional
rlabel 
 s 0 15 24 18 6 VDDA
port 5 nsew power bidirectional
rlabel 
 s 50 15 74 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 15 24 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 50 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 17 74 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 17 74 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 17 74 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 17 74 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 17 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 17 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 17 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 17 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 18 73 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 18 73 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 17 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 17 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 73 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 17 72 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 17 72 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 17 72 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 17 72 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 17 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 17 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 17 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 17 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 18 71 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 18 71 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 17 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 17 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 71 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 17 70 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 17 70 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 17 70 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 17 70 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 17 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 17 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 17 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 17 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 18 69 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 18 69 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 17 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 17 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 69 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 17 68 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 17 68 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 17 68 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 17 68 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 17 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 17 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 17 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 17 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 18 67 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 18 67 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 17 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 17 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 67 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 18 66 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 18 66 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 17 66 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 17 66 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 66 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 18 66 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 18 66 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 17 66 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 17 66 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 66 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 17 65 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 17 65 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 17 65 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 17 65 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 17 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 17 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 17 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 17 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 18 64 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 18 64 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 17 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 17 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 64 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 17 63 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 17 63 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 17 63 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 17 63 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 17 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 17 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 17 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 17 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 18 62 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 18 62 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 17 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 17 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 62 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 17 61 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 17 61 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 17 61 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 17 61 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 17 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 17 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 17 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 17 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 18 60 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 18 60 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 17 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 17 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 60 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 17 59 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 17 59 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 17 59 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 17 59 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 17 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 17 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 17 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 17 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 18 58 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 18 58 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 17 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 17 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 58 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 17 57 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 17 57 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 17 57 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 17 57 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 17 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 17 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 17 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 17 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 18 56 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 18 56 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 17 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 17 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 56 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 18 55 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 18 55 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 17 55 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 17 55 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 18 55 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 18 55 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 17 55 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 17 55 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 17 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 17 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 17 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 17 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 18 54 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 18 54 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 17 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 17 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 54 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 17 53 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 17 53 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 53 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 17 53 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 17 53 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 53 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 17 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 17 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 17 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 17 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 18 52 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 18 52 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 17 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 17 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 52 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 18 51 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 18 51 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 17 51 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 17 51 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 51 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 18 51 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 18 51 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 17 51 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 17 51 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 16 51 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 16 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 15 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 50 15 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 17 24 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 17 24 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 17 24 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 17 24 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 17 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 17 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 17 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 17 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 18 23 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 18 23 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 17 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 17 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 23 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 17 22 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 17 22 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 17 22 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 17 22 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 17 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 17 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 17 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 17 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 18 21 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 18 21 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 17 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 17 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 21 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 17 20 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 17 20 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 17 20 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 17 20 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 17 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 17 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 17 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 17 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 18 19 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 18 19 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 17 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 17 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 19 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 17 18 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 17 18 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 17 18 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 17 18 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 17 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 17 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 17 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 17 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 18 17 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 18 17 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 17 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 17 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 17 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 17 16 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 17 16 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 17 16 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 17 16 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 17 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 17 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 17 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 17 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 18 15 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 18 15 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 17 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 17 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 15 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 17 14 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 17 14 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 17 14 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 17 14 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 17 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 17 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 17 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 17 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 18 13 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 18 13 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 17 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 17 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 13 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 17 12 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 17 12 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 17 12 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 17 12 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 17 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 17 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 17 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 17 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 18 11 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 18 11 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 17 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 17 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 11 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 17 10 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 17 10 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 17 10 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 17 10 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 17 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 17 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 17 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 17 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 18 9 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 18 9 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 17 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 17 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 9 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 17 8 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 17 8 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 17 8 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 17 8 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 17 7 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 17 7 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 17 7 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 17 7 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 17 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 17 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 17 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 17 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 18 6 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 18 6 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 17 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 17 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 6 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 17 5 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 17 5 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 17 5 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 17 5 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 17 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 17 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 17 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 17 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 18 4 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 18 4 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 17 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 17 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 4 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 17 3 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 17 3 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 17 3 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 17 3 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 17 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 17 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 17 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 17 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 18 2 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 18 2 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 17 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 17 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 2 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 17 1 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 17 1 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 17 1 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 17 1 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 17 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 69 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 64 1 68 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 64 75 68 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 1 48 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 52 1 53 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 56 1 57 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 48 75 48 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 52 75 53 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 56 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 48 1 57 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 48 75 57 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 200
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
