magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 30 43 764 283
rect -26 -43 794 43
<< locali >>
rect 208 420 274 751
rect 536 420 586 751
rect 208 386 743 420
rect 25 316 567 350
rect 603 310 743 386
rect 603 280 637 310
rect 208 246 637 280
rect 208 99 258 246
rect 520 99 637 246
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 18 735 136 751
rect 18 701 24 735
rect 58 701 96 735
rect 130 701 136 735
rect 18 435 136 701
rect 310 735 500 751
rect 310 701 316 735
rect 350 701 388 735
rect 422 701 460 735
rect 494 701 500 735
rect 310 456 500 701
rect 624 735 742 751
rect 624 701 630 735
rect 664 701 702 735
rect 736 701 742 735
rect 624 456 742 701
rect 18 113 136 265
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 136 113
rect 294 113 484 210
rect 18 73 136 79
rect 294 79 300 113
rect 334 79 372 113
rect 406 79 444 113
rect 478 79 484 113
rect 676 113 742 265
rect 294 73 484 79
rect 676 79 682 113
rect 716 79 742 113
rect 676 73 742 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 24 701 58 735
rect 96 701 130 735
rect 316 701 350 735
rect 388 701 422 735
rect 460 701 494 735
rect 630 701 664 735
rect 702 701 736 735
rect 24 79 58 113
rect 96 79 130 113
rect 300 79 334 113
rect 372 79 406 113
rect 444 79 478 113
rect 682 79 716 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 316 735
rect 350 701 388 735
rect 422 701 460 735
rect 494 701 630 735
rect 664 701 702 735
rect 736 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 300 113
rect 334 79 372 113
rect 406 79 444 113
rect 478 79 682 113
rect 716 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel locali s 25 316 567 350 6 A
port 1 nsew signal input
rlabel metal1 s 0 51 768 125 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 768 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 794 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 30 43 764 283 6 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 768 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 834 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 768 763 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 520 99 637 246 6 Y
port 6 nsew signal output
rlabel locali s 208 99 258 246 6 Y
port 6 nsew signal output
rlabel locali s 208 246 637 280 6 Y
port 6 nsew signal output
rlabel locali s 603 280 637 310 6 Y
port 6 nsew signal output
rlabel locali s 603 310 743 386 6 Y
port 6 nsew signal output
rlabel locali s 208 386 743 420 6 Y
port 6 nsew signal output
rlabel locali s 536 420 586 751 6 Y
port 6 nsew signal output
rlabel locali s 208 420 274 751 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 768 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 69816
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 59660
<< end >>
