magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 3 11 6 6 DRAIN
port 1 nsew
rlabel  s 2 8 10 9 6 GATE
port 2 nsew
rlabel  s 2 0 10 1 8 GATE
port 2 nsew
rlabel  s 0 6 11 8 6 SOURCE
port 3 nsew
rlabel  s 0 1 11 3 6 SOURCE
port 3 nsew
rlabel  s 0 1 1 8 4 SUBSTRATE
port 4 nsew
rlabel  s 11 1 11 8 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 11 9
string LEFview TRUE
<< end >>
