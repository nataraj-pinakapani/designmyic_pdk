magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< poly >>
rect -13 6277 147 6293
rect -13 6243 16 6277
rect 50 6243 84 6277
rect 118 6243 147 6277
rect -13 3809 16 3843
rect 50 3809 84 3843
rect 118 3809 147 3843
rect -13 3793 147 3809
rect 278 6180 438 6196
rect 278 6146 307 6180
rect 341 6146 375 6180
rect 409 6146 438 6180
rect -13 3705 147 3721
rect -13 3671 16 3705
rect 50 3671 84 3705
rect 118 3671 147 3705
rect -283 3416 -123 3432
rect -283 3382 -254 3416
rect -220 3382 -186 3416
rect -152 3382 -123 3416
rect -283 3048 -254 3082
rect -220 3048 -186 3082
rect -152 3048 -123 3082
rect -283 3032 -123 3048
rect -283 2831 -123 2847
rect -283 2797 -254 2831
rect -220 2797 -186 2831
rect -152 2797 -123 2831
rect -283 2463 -254 2497
rect -220 2463 -186 2497
rect -152 2463 -123 2497
rect -283 2447 -123 2463
rect -13 2437 16 2471
rect 50 2437 84 2471
rect 118 2437 147 2471
rect -13 2421 147 2437
rect -13 2363 147 2379
rect -13 2329 16 2363
rect 50 2329 84 2363
rect 118 2329 147 2363
rect -281 2275 -121 2291
rect -281 2241 -252 2275
rect -218 2241 -184 2275
rect -150 2241 -121 2275
rect -281 1907 -252 1941
rect -218 1907 -184 1941
rect -150 1907 -121 1941
rect -281 1891 -121 1907
rect -281 1690 -121 1706
rect -281 1656 -252 1690
rect -218 1656 -184 1690
rect -150 1656 -121 1690
rect -281 1322 -252 1356
rect -218 1322 -184 1356
rect -150 1322 -121 1356
rect -281 1306 -121 1322
rect -13 1095 16 1129
rect 50 1095 84 1129
rect 118 1095 147 1129
rect 534 6180 694 6196
rect 534 6146 563 6180
rect 597 6146 631 6180
rect 665 6146 694 6180
rect -13 1079 147 1095
<< polycont >>
rect 16 6243 50 6277
rect 84 6243 118 6277
rect 16 3809 50 3843
rect 84 3809 118 3843
rect 307 6146 341 6180
rect 375 6146 409 6180
rect 16 3671 50 3705
rect 84 3671 118 3705
rect -254 3382 -220 3416
rect -186 3382 -152 3416
rect -254 3048 -220 3082
rect -186 3048 -152 3082
rect -254 2797 -220 2831
rect -186 2797 -152 2831
rect -254 2463 -220 2497
rect -186 2463 -152 2497
rect 16 2437 50 2471
rect 84 2437 118 2471
rect 16 2329 50 2363
rect 84 2329 118 2363
rect -252 2241 -218 2275
rect -184 2241 -150 2275
rect -252 1907 -218 1941
rect -184 1907 -150 1941
rect -252 1656 -218 1690
rect -184 1656 -150 1690
rect -252 1322 -218 1356
rect -184 1322 -150 1356
rect 16 1095 50 1129
rect 84 1095 118 1129
rect 563 6146 597 6180
rect 631 6146 665 6180
<< npolyres >>
rect -13 3843 147 6243
rect -283 3082 -123 3382
rect -283 2497 -123 2797
rect -13 2471 147 3671
rect -281 1941 -121 2241
rect -281 1356 -121 1656
rect -13 1129 147 2329
rect 278 1274 438 6146
rect 534 1274 694 6146
rect 278 1114 694 1274
<< locali >>
rect -1 6277 425 6278
rect -1 6243 16 6277
rect 50 6271 84 6277
rect 118 6271 425 6277
rect -1 6093 17 6243
rect 411 6093 425 6271
rect 547 6146 563 6180
rect 597 6146 631 6180
rect 665 6146 681 6180
rect -1 5670 425 6093
rect 0 3677 14 3843
rect 120 3677 134 3843
rect 0 3671 16 3677
rect 50 3671 84 3677
rect 118 3671 134 3677
rect -270 3382 -254 3588
rect -148 3410 -136 3588
rect -220 3382 -186 3410
rect -152 3382 -136 3410
rect -270 3048 -256 3082
rect -220 3048 -186 3082
rect -150 3048 -136 3082
rect -270 2964 -136 3048
rect -270 2858 -256 2964
rect -150 2858 -136 2964
rect -270 2831 -136 2858
rect -270 2797 -254 2831
rect -220 2797 -186 2831
rect -152 2797 -136 2831
rect -270 2463 -256 2497
rect -220 2463 -186 2497
rect -150 2463 -136 2497
rect -270 2275 -136 2463
rect 0 2437 14 2471
rect 120 2437 134 2471
rect 0 2363 131 2437
rect 0 2329 14 2363
rect 50 2329 84 2363
rect 120 2329 134 2363
rect -270 2241 -254 2275
rect -218 2241 -184 2275
rect -148 2241 -134 2275
rect -268 1911 -252 1941
rect -218 1911 -184 1941
rect -150 1911 -134 1941
rect -268 1805 -254 1911
rect -148 1805 -134 1911
rect -268 1711 -134 1805
rect -268 1677 -254 1711
rect -220 1690 -182 1711
rect -268 1656 -252 1677
rect -218 1656 -184 1690
rect -148 1677 -134 1711
rect -150 1656 -134 1677
rect -268 1349 -252 1356
rect -218 1349 -184 1356
rect -268 1243 -256 1349
rect -150 1243 -134 1356
rect 0 1273 134 1279
rect 0 1095 14 1273
rect 120 1095 134 1273
<< viali >>
rect 17 6243 50 6271
rect 50 6243 84 6271
rect 84 6243 118 6271
rect 118 6243 411 6271
rect 17 6180 411 6243
rect 17 6146 307 6180
rect 307 6146 341 6180
rect 341 6146 375 6180
rect 375 6146 409 6180
rect 409 6146 411 6180
rect 17 6093 411 6146
rect 14 3843 120 3855
rect 14 3809 16 3843
rect 16 3809 50 3843
rect 50 3809 84 3843
rect 84 3809 118 3843
rect 118 3809 120 3843
rect 14 3705 120 3809
rect 14 3677 16 3705
rect 16 3677 50 3705
rect 50 3677 84 3705
rect 84 3677 118 3705
rect 118 3677 120 3705
rect -254 3416 -148 3588
rect -254 3410 -220 3416
rect -220 3410 -186 3416
rect -186 3410 -152 3416
rect -152 3410 -148 3416
rect -256 3048 -254 3082
rect -254 3048 -222 3082
rect -184 3048 -152 3082
rect -152 3048 -150 3082
rect -256 2858 -150 2964
rect -256 2463 -254 2497
rect -254 2463 -222 2497
rect -184 2463 -152 2497
rect -152 2463 -150 2497
rect 14 2471 120 2615
rect 14 2437 16 2471
rect 16 2437 50 2471
rect 50 2437 84 2471
rect 84 2437 118 2471
rect 118 2437 120 2471
rect 14 2329 16 2363
rect 16 2329 48 2363
rect 86 2329 118 2363
rect 118 2329 120 2363
rect -254 2241 -252 2275
rect -252 2241 -220 2275
rect -182 2241 -150 2275
rect -150 2241 -148 2275
rect -254 1907 -252 1911
rect -252 1907 -218 1911
rect -218 1907 -184 1911
rect -184 1907 -150 1911
rect -150 1907 -148 1911
rect -254 1805 -148 1907
rect -254 1690 -220 1711
rect -182 1690 -148 1711
rect -254 1677 -252 1690
rect -252 1677 -220 1690
rect -182 1677 -150 1690
rect -150 1677 -148 1690
rect -256 1322 -252 1349
rect -252 1322 -218 1349
rect -218 1322 -184 1349
rect -184 1322 -150 1349
rect -256 1171 -150 1322
rect 14 1129 120 1273
rect 14 1095 16 1129
rect 16 1095 50 1129
rect 50 1095 84 1129
rect 84 1095 118 1129
rect 118 1095 120 1129
<< metal1 >>
rect 5 6271 423 6277
rect 5 6093 17 6271
rect 411 6093 423 6271
rect 5 6087 423 6093
rect 2 3855 132 3861
rect 2 3677 14 3855
rect 120 3677 132 3855
rect 2 3619 132 3677
rect 3 3617 131 3618
rect -268 3564 -262 3616
rect -210 3588 -194 3616
rect -142 3564 -136 3616
rect -268 3546 -254 3564
rect -148 3546 -136 3564
rect -268 3494 -262 3546
rect -142 3494 -136 3546
rect -268 3410 -254 3494
rect -148 3410 -136 3494
rect -268 3396 -136 3410
rect -267 3394 -137 3395
rect -268 3094 -136 3394
rect -267 3093 -137 3094
rect -268 3082 -136 3092
rect -268 3048 -256 3082
rect -222 3048 -184 3082
rect -150 3048 -136 3082
rect -268 2964 -136 3048
rect -268 2858 -256 2964
rect -150 2858 -136 2964
rect -268 2815 -136 2858
rect -267 2813 -137 2814
rect -268 2513 -136 2813
rect -267 2512 -137 2513
rect -268 2497 -136 2511
rect -268 2463 -256 2497
rect -222 2463 -184 2497
rect -150 2463 -136 2497
rect -268 2275 -136 2463
rect -268 2241 -254 2275
rect -220 2241 -182 2275
rect -148 2241 -136 2275
rect -268 2226 -136 2241
rect -267 2224 -137 2225
rect -268 1924 -136 2224
rect -267 1923 -137 1924
rect -268 1911 -136 1922
rect -268 1805 -254 1911
rect -148 1805 -136 1911
rect -268 1711 -136 1805
rect -268 1677 -254 1711
rect -220 1677 -182 1711
rect -148 1677 -136 1711
rect -268 1666 -136 1677
rect -267 1664 -137 1665
rect -268 1364 -136 1664
rect -267 1363 -137 1364
rect -268 1349 -136 1362
rect -268 1171 -256 1349
rect -150 1310 -136 1349
rect 3 3580 131 3581
rect 2 2615 132 3579
rect 2 2437 14 2615
rect 120 2437 132 2615
rect 2 2363 132 2437
rect 2 2329 14 2363
rect 48 2329 86 2363
rect 120 2329 132 2363
rect 2 2271 132 2329
rect 3 2269 131 2270
rect 2 2233 132 2269
rect 3 2232 131 2233
rect 2 2133 132 2231
rect 2 2081 8 2133
rect 60 2081 74 2133
rect 126 2081 132 2133
rect 2 2063 132 2081
rect 2 2011 8 2063
rect 60 2011 74 2063
rect 126 2011 132 2063
rect 209 3564 215 3616
rect 267 3564 285 3616
rect 209 3546 285 3564
rect 209 3494 215 3546
rect 267 3494 285 3546
rect 209 2133 285 3494
rect 209 2081 215 2133
rect 267 2081 285 2133
rect 209 2063 285 2081
rect 209 2011 215 2063
rect 267 2011 285 2063
rect -150 1171 -138 1310
rect -268 1165 -138 1171
rect 2 1273 132 2011
rect 2 1095 14 1273
rect 120 1095 132 1273
rect 2 1089 132 1095
<< rmetal1 >>
rect 2 3618 132 3619
rect 2 3617 3 3618
rect 131 3617 132 3618
rect -268 3395 -136 3396
rect -268 3394 -267 3395
rect -137 3394 -136 3395
rect -268 3093 -267 3094
rect -137 3093 -136 3094
rect -268 3092 -136 3093
rect -268 2814 -136 2815
rect -268 2813 -267 2814
rect -137 2813 -136 2814
rect -268 2512 -267 2513
rect -137 2512 -136 2513
rect -268 2511 -136 2512
rect -268 2225 -136 2226
rect -268 2224 -267 2225
rect -137 2224 -136 2225
rect -268 1923 -267 1924
rect -137 1923 -136 1924
rect -268 1922 -136 1923
rect -268 1665 -136 1666
rect -268 1664 -267 1665
rect -137 1664 -136 1665
rect -268 1363 -267 1364
rect -137 1363 -136 1364
rect -268 1362 -136 1363
rect 2 3580 3 3581
rect 131 3580 132 3581
rect 2 3579 132 3580
rect 2 2270 132 2271
rect 2 2269 3 2270
rect 131 2269 132 2270
rect 2 2232 3 2233
rect 131 2232 132 2233
rect 2 2231 132 2232
<< via1 >>
rect -262 3588 -210 3616
rect -194 3588 -142 3616
rect -262 3564 -254 3588
rect -254 3564 -210 3588
rect -194 3564 -148 3588
rect -148 3564 -142 3588
rect -262 3494 -254 3546
rect -254 3494 -210 3546
rect -194 3494 -148 3546
rect -148 3494 -142 3546
rect 8 2081 60 2133
rect 74 2081 126 2133
rect 8 2011 60 2063
rect 74 2011 126 2063
rect 215 3564 267 3616
rect 215 3494 267 3546
rect 215 2081 267 2133
rect 215 2011 267 2063
<< metal2 >>
rect -268 3564 -262 3616
rect -210 3564 -194 3616
rect -142 3564 215 3616
rect 267 3564 285 3616
rect -268 3546 285 3564
rect -268 3494 -262 3546
rect -210 3494 -194 3546
rect -142 3494 215 3546
rect 267 3494 285 3546
rect 2 2081 8 2133
rect 60 2081 74 2133
rect 126 2081 215 2133
rect 267 2081 285 2133
rect 2 2063 285 2081
rect 2 2011 8 2063
rect 60 2011 74 2063
rect 126 2011 215 2063
rect 267 2011 285 2063
use sky130_fd_io__tk_em1o_cdns_55959141808289  sky130_fd_io__tk_em1o_cdns_55959141808289_0
timestamp 1663361622
transform 0 1 2 -1 0 3671
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_0
timestamp 1663361622
transform 0 1 -268 -1 0 3448
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_1
timestamp 1663361622
transform 0 1 -268 -1 0 2867
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_2
timestamp 1663361622
transform 0 -1 -136 -1 0 1718
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_3
timestamp 1663361622
transform 0 -1 -136 -1 0 2278
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_0
timestamp 1663361622
transform 0 1 2 -1 0 2323
box 0 0 1 1
use sky130_fd_pr__res_bent_po__example_5595914180862  sky130_fd_pr__res_bent_po__example_5595914180862_0
timestamp 1663361622
transform 0 1 -13 -1 0 2329
box -50 13 1185 14
use sky130_fd_pr__res_bent_po__example_5595914180862  sky130_fd_pr__res_bent_po__example_5595914180862_1
timestamp 1663361622
transform 0 1 -13 -1 0 3671
box -50 13 1185 14
use sky130_fd_pr__res_bent_po__example_5595914180863  sky130_fd_pr__res_bent_po__example_5595914180863_0
timestamp 1663361622
transform 0 -1 147 1 0 3843
box -50 13 2385 14
use sky130_fd_pr__res_bent_po__example_55959141808715  sky130_fd_pr__res_bent_po__example_55959141808715_0
timestamp 1663361622
transform 0 -1 438 -1 0 6146
box -50 -243 -49 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_0
timestamp 1663361622
transform 0 1 -283 -1 0 3382
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_1
timestamp 1663361622
transform 0 1 -283 -1 0 2797
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_2
timestamp 1663361622
transform 0 -1 -121 -1 0 1656
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_3
timestamp 1663361622
transform 0 -1 -121 -1 0 2241
box 15 13 285 14
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1663361622
transform 1 0 -256 0 1 3048
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1663361622
transform 1 0 -256 0 1 2463
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1663361622
transform -1 0 -148 0 1 1677
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1663361622
transform -1 0 -148 0 -1 2275
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1663361622
transform 1 0 -256 0 1 2858
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_1
timestamp 1663361622
transform -1 0 -148 0 -1 1911
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_0
timestamp 1663361622
transform -1 0 120 0 -1 1273
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_1
timestamp 1663361622
transform 1 0 -254 0 1 3410
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_2
timestamp 1663361622
transform -1 0 -150 0 1 1171
box 0 0 1 1
<< labels >>
<< properties >>
string GDS_END 3929200
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 3921810
<< end >>
