magic
tech sky130A
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__dfm1sd__example_55959141808258  sky130_fd_pr__dfm1sd__example_55959141808258_0
timestamp 1663361622
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180893  sky130_fd_pr__hvdfm1sd__example_5595914180893_0
timestamp 1663361622
transform 1 0 1600 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 32707088
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 32706164
<< end >>
