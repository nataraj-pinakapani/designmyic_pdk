magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 1 0 2 4 6 C0
port 1 nsew
rlabel  s 1 0 1 4 6 C0
port 1 nsew
rlabel  s 0 0 0 4 4 C0
port 1 nsew
rlabel  s 0 0 2 0 8 C0
port 1 nsew
rlabel  s 2 0 2 4 6 C1
port 2 nsew
rlabel  s 1 0 1 4 6 C1
port 2 nsew
rlabel  s 1 0 1 4 6 C1
port 2 nsew
rlabel  s 0 0 0 4 4 C1
port 2 nsew
rlabel  s 0 4 2 5 6 C1
port 2 nsew
rlabel  s 0 0 0 4 4 C1
port 2 nsew
rlabel metal_blue s 0 2 1 3 4 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 2 5
string LEFview TRUE
<< end >>
