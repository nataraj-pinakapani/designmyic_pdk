magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< locali >>
rect 12165 1381 12231 1473
rect 12178 1347 12216 1381
<< viali >>
rect 12144 1347 12178 1381
rect 12216 1347 12250 1381
<< metal1 >>
rect 2787 2731 3539 2732
rect 2787 2679 2793 2731
rect 2845 2679 2892 2731
rect 2944 2679 2991 2731
rect 3043 2679 3089 2731
rect 3141 2679 3187 2731
rect 3239 2679 3285 2731
rect 3337 2679 3383 2731
rect 3435 2679 3481 2731
rect 3533 2679 3539 2731
rect 2787 2643 3539 2679
rect 2787 2591 2793 2643
rect 2845 2591 2892 2643
rect 2944 2591 2991 2643
rect 3043 2591 3089 2643
rect 3141 2591 3187 2643
rect 3239 2591 3285 2643
rect 3337 2591 3383 2643
rect 3435 2591 3481 2643
rect 3533 2591 3539 2643
rect 2787 2555 3539 2591
rect 5273 2579 5506 2710
rect 2787 2503 2793 2555
rect 2845 2503 2892 2555
rect 2944 2503 2991 2555
rect 3043 2503 3089 2555
rect 3141 2503 3187 2555
rect 3239 2503 3285 2555
rect 3337 2503 3383 2555
rect 3435 2503 3481 2555
rect 3533 2503 3539 2555
rect 2787 2502 3539 2503
rect 11522 2498 11542 2700
rect 12400 2498 12458 2700
rect 14371 2498 14400 2700
rect 11522 2424 11542 2470
rect 12400 2424 12458 2470
rect 14371 2424 14400 2470
rect 3224 2201 3334 2247
rect 3689 2037 3741 2043
rect 3689 1973 3741 1985
rect 2858 1906 2864 1958
rect 2916 1906 2928 1958
rect 2980 1906 2986 1958
rect 3122 1905 3128 1957
rect 3180 1905 3198 1957
rect 3250 1905 3267 1957
rect 3319 1905 3336 1957
rect 3388 1905 3394 1957
rect 11555 1972 11581 2248
rect 12400 1972 12429 2248
rect 14371 1972 14400 2248
tri 3687 1915 3689 1917 se
rect 3689 1915 3741 1921
tri 3678 1906 3687 1915 se
rect 3687 1906 3741 1915
rect 3879 1906 3885 1958
rect 3937 1906 3949 1958
rect 4001 1906 4007 1958
tri 3677 1905 3678 1906 se
rect 3678 1905 3741 1906
tri 3667 1895 3677 1905 se
rect 3677 1895 3741 1905
tri 3638 1866 3667 1895 se
rect 3667 1880 3726 1895
tri 3726 1880 3741 1895 nw
rect 4887 1880 4893 1932
rect 4945 1880 4957 1932
rect 5009 1880 5015 1932
rect 11142 1904 12092 1944
rect 3667 1871 3717 1880
tri 3717 1871 3726 1880 nw
rect 3667 1866 3712 1871
tri 3712 1866 3717 1871 nw
rect 3236 1814 3242 1866
rect 3294 1814 3306 1866
rect 3358 1843 3689 1866
tri 3689 1843 3712 1866 nw
rect 3358 1821 3667 1843
tri 3667 1821 3689 1843 nw
rect 10588 1821 10594 1873
rect 10646 1821 10658 1873
rect 10710 1821 10716 1873
rect 10843 1821 10849 1873
rect 10901 1821 10913 1873
rect 10965 1821 10971 1873
rect 3358 1814 3660 1821
tri 3660 1814 3667 1821 nw
rect 7703 1643 7781 1749
rect 10633 1720 10685 1821
rect 10578 1668 10584 1720
rect 10636 1668 10648 1720
rect 10700 1668 10706 1720
rect 10843 1707 10971 1821
rect 2773 1578 2779 1630
rect 2831 1578 2864 1630
rect 2916 1578 2949 1630
rect 3001 1578 3007 1630
rect 2773 1558 3007 1578
rect 2773 1506 2779 1558
rect 2831 1506 2864 1558
rect 2916 1506 2949 1558
rect 3001 1506 3007 1558
rect 3061 1511 3294 1626
rect 7685 1591 7691 1643
rect 7743 1591 7755 1643
rect 7807 1591 7813 1643
rect 10843 1639 10942 1707
tri 10942 1678 10971 1707 nw
rect 4449 1500 4455 1552
rect 4507 1500 4525 1552
rect 4577 1500 4595 1552
rect 4647 1500 4665 1552
rect 4717 1500 4735 1552
rect 4787 1500 4805 1552
rect 4857 1500 4875 1552
rect 4927 1500 4944 1552
rect 4996 1500 5002 1552
rect 8613 1547 8663 1593
rect 10814 1587 10820 1639
rect 10872 1587 10884 1639
rect 10936 1587 10942 1639
rect 5354 1505 5412 1547
rect 10820 1452 10872 1458
rect 11142 1427 11182 1904
rect 10872 1400 11182 1427
rect 10820 1388 11182 1400
rect 10872 1387 11182 1388
rect 11248 1837 11300 1843
rect 13410 1819 13416 1871
rect 13468 1819 13480 1871
rect 13532 1819 13538 1871
rect 11248 1773 11300 1785
rect 13467 1734 13473 1786
rect 13525 1734 13537 1786
rect 13589 1734 13595 1786
rect 11248 1387 11300 1721
rect 13467 1654 13473 1706
rect 13525 1654 13537 1706
rect 13589 1654 13595 1706
rect 14219 1574 14225 1626
rect 14277 1574 14289 1626
rect 14341 1574 14347 1626
rect 12939 1520 12978 1541
rect 12679 1475 12721 1503
rect 12911 1492 13039 1520
rect 14236 1415 14338 1447
rect 11248 1381 12262 1387
rect 11248 1354 12144 1381
rect 12132 1347 12144 1354
rect 12178 1347 12216 1381
rect 12250 1347 12262 1381
rect 12132 1341 12262 1347
rect 10820 1330 10872 1336
rect 9612 1287 9670 1329
rect 4800 823 5019 1016
<< via1 >>
rect 2793 2679 2845 2731
rect 2892 2679 2944 2731
rect 2991 2679 3043 2731
rect 3089 2679 3141 2731
rect 3187 2679 3239 2731
rect 3285 2679 3337 2731
rect 3383 2679 3435 2731
rect 3481 2679 3533 2731
rect 2793 2591 2845 2643
rect 2892 2591 2944 2643
rect 2991 2591 3043 2643
rect 3089 2591 3141 2643
rect 3187 2591 3239 2643
rect 3285 2591 3337 2643
rect 3383 2591 3435 2643
rect 3481 2591 3533 2643
rect 2793 2503 2845 2555
rect 2892 2503 2944 2555
rect 2991 2503 3043 2555
rect 3089 2503 3141 2555
rect 3187 2503 3239 2555
rect 3285 2503 3337 2555
rect 3383 2503 3435 2555
rect 3481 2503 3533 2555
rect 3689 1985 3741 2037
rect 2864 1906 2916 1958
rect 2928 1906 2980 1958
rect 3128 1905 3180 1957
rect 3198 1905 3250 1957
rect 3267 1905 3319 1957
rect 3336 1905 3388 1957
rect 3689 1921 3741 1973
rect 3885 1906 3937 1958
rect 3949 1906 4001 1958
rect 4893 1880 4945 1932
rect 4957 1880 5009 1932
rect 3242 1814 3294 1866
rect 3306 1814 3358 1866
rect 10594 1821 10646 1873
rect 10658 1821 10710 1873
rect 10849 1821 10901 1873
rect 10913 1821 10965 1873
rect 10584 1668 10636 1720
rect 10648 1668 10700 1720
rect 2779 1578 2831 1630
rect 2864 1578 2916 1630
rect 2949 1578 3001 1630
rect 2779 1506 2831 1558
rect 2864 1506 2916 1558
rect 2949 1506 3001 1558
rect 7691 1591 7743 1643
rect 7755 1591 7807 1643
rect 4455 1500 4507 1552
rect 4525 1500 4577 1552
rect 4595 1500 4647 1552
rect 4665 1500 4717 1552
rect 4735 1500 4787 1552
rect 4805 1500 4857 1552
rect 4875 1500 4927 1552
rect 4944 1500 4996 1552
rect 10820 1587 10872 1639
rect 10884 1587 10936 1639
rect 10820 1400 10872 1452
rect 10820 1336 10872 1388
rect 11248 1785 11300 1837
rect 13416 1819 13468 1871
rect 13480 1819 13532 1871
rect 11248 1721 11300 1773
rect 13473 1734 13525 1786
rect 13537 1734 13589 1786
rect 13473 1654 13525 1706
rect 13537 1654 13589 1706
rect 14225 1574 14277 1626
rect 14289 1574 14341 1626
<< metal2 >>
rect 2779 2676 2788 2732
rect 2844 2731 2874 2732
rect 2930 2731 2960 2732
rect 3016 2731 3046 2732
rect 3102 2731 3131 2732
rect 3187 2731 3216 2732
rect 3272 2731 3301 2732
rect 3357 2731 3386 2732
rect 2845 2679 2874 2731
rect 2944 2679 2960 2731
rect 3043 2679 3046 2731
rect 3272 2679 3285 2731
rect 3357 2679 3383 2731
rect 2844 2676 2874 2679
rect 2930 2676 2960 2679
rect 3016 2676 3046 2679
rect 3102 2676 3131 2679
rect 3187 2676 3216 2679
rect 3272 2676 3301 2679
rect 3357 2676 3386 2679
rect 3442 2676 3471 2732
rect 3527 2731 3539 2732
rect 3533 2679 3539 2731
rect 3527 2676 3539 2679
rect 2779 2648 3539 2676
rect 2779 2592 2788 2648
rect 2844 2643 2874 2648
rect 2930 2643 2960 2648
rect 3016 2643 3046 2648
rect 3102 2643 3131 2648
rect 3187 2643 3216 2648
rect 3272 2643 3301 2648
rect 3357 2643 3386 2648
rect 2845 2592 2874 2643
rect 2944 2592 2960 2643
rect 3043 2592 3046 2643
rect 3272 2592 3285 2643
rect 3357 2592 3383 2643
rect 3442 2592 3471 2648
rect 3527 2643 3539 2648
rect 2779 2591 2793 2592
rect 2845 2591 2892 2592
rect 2944 2591 2991 2592
rect 3043 2591 3089 2592
rect 3141 2591 3187 2592
rect 3239 2591 3285 2592
rect 3337 2591 3383 2592
rect 3435 2591 3481 2592
rect 3533 2591 3539 2643
rect 2779 2564 3539 2591
rect 2779 2508 2788 2564
rect 2844 2555 2874 2564
rect 2930 2555 2960 2564
rect 3016 2555 3046 2564
rect 3102 2555 3131 2564
rect 3187 2555 3216 2564
rect 3272 2555 3301 2564
rect 3357 2555 3386 2564
rect 2845 2508 2874 2555
rect 2944 2508 2960 2555
rect 3043 2508 3046 2555
rect 3272 2508 3285 2555
rect 3357 2508 3383 2555
rect 3442 2508 3471 2564
rect 3527 2555 3539 2564
rect 2787 2503 2793 2508
rect 2845 2503 2892 2508
rect 2944 2503 2991 2508
rect 3043 2503 3089 2508
rect 3141 2503 3187 2508
rect 3239 2503 3285 2508
rect 3337 2503 3383 2508
rect 3435 2503 3481 2508
rect 3533 2503 3539 2555
rect 2787 2502 3539 2503
tri 3007 2041 3010 2044 se
rect 3010 2041 3518 2044
tri 3518 2041 3521 2044 sw
tri 3003 2037 3007 2041 se
rect 3007 2037 3521 2041
tri 3521 2037 3525 2041 sw
rect 3689 2040 4181 2073
tri 4181 2040 4214 2073 sw
rect 3689 2037 6615 2040
tri 2951 1985 3003 2037 se
rect 3003 2004 3525 2037
rect 3003 1985 3037 2004
tri 3037 1985 3056 2004 nw
tri 3476 1985 3495 2004 ne
rect 3495 1985 3525 2004
tri 3525 1985 3577 2037 sw
rect 3741 2031 6615 2037
tri 4165 1998 4198 2031 ne
rect 4198 2002 6615 2031
tri 6615 2002 6653 2040 sw
rect 4198 1998 6653 2002
tri 2939 1973 2951 1985 se
rect 2951 1973 3025 1985
tri 3025 1973 3037 1985 nw
tri 3495 1973 3507 1985 ne
rect 3507 1973 3577 1985
tri 3577 1973 3589 1985 sw
rect 3689 1973 3741 1985
tri 2925 1959 2939 1973 se
rect 2939 1959 3011 1973
tri 3011 1959 3025 1973 nw
tri 3507 1959 3521 1973 ne
rect 3521 1959 3589 1973
tri 3589 1959 3603 1973 sw
tri 2924 1958 2925 1959 se
rect 2925 1958 3010 1959
tri 3010 1958 3011 1959 nw
tri 3521 1958 3522 1959 ne
rect 3522 1958 3603 1959
tri 3603 1958 3604 1959 sw
rect 2858 1906 2864 1958
rect 2916 1906 2928 1958
rect 2980 1957 3009 1958
tri 3009 1957 3010 1958 nw
tri 3522 1957 3523 1958 ne
rect 3523 1957 3604 1958
tri 3604 1957 3605 1958 sw
rect 2980 1906 2986 1957
tri 2986 1934 3009 1957 nw
rect 3122 1905 3128 1957
rect 3180 1905 3198 1957
rect 3250 1905 3267 1957
rect 3319 1905 3336 1957
rect 3388 1934 3471 1957
tri 3471 1934 3494 1957 sw
tri 3523 1934 3546 1957 ne
rect 3546 1934 3605 1957
rect 3388 1928 3494 1934
tri 3494 1928 3500 1934 sw
tri 3546 1928 3552 1934 ne
rect 3552 1928 3605 1934
rect 3388 1921 3500 1928
tri 3500 1921 3507 1928 sw
tri 3552 1921 3559 1928 ne
rect 3559 1921 3605 1928
tri 3605 1921 3641 1957 sw
tri 6599 1958 6639 1998 ne
rect 6639 1958 6653 1998
rect 3388 1906 3507 1921
tri 3507 1906 3522 1921 sw
tri 3559 1906 3574 1921 ne
rect 3574 1915 3641 1921
tri 3641 1915 3647 1921 sw
rect 3689 1915 3741 1921
rect 3574 1906 3647 1915
tri 3647 1906 3656 1915 sw
rect 3879 1906 3885 1958
rect 3937 1906 3949 1958
rect 4001 1906 4007 1958
tri 6639 1944 6653 1958 ne
tri 6653 1944 6711 2002 sw
tri 6653 1932 6665 1944 ne
rect 6665 1932 11181 1944
rect 3388 1905 3522 1906
tri 3522 1905 3523 1906 sw
tri 3574 1905 3575 1906 ne
rect 3575 1905 3656 1906
tri 3656 1905 3657 1906 sw
tri 3465 1880 3490 1905 ne
rect 3490 1880 3523 1905
tri 3523 1880 3548 1905 sw
tri 3575 1880 3600 1905 ne
rect 3600 1880 3657 1905
tri 3657 1880 3682 1905 sw
tri 3490 1876 3494 1880 ne
rect 3494 1877 3548 1880
tri 3548 1877 3551 1880 sw
tri 3600 1877 3603 1880 ne
rect 3603 1877 3682 1880
tri 3682 1877 3685 1880 sw
rect 3494 1876 3551 1877
tri 3551 1876 3552 1877 sw
tri 3603 1876 3604 1877 ne
rect 3604 1876 3685 1877
tri 3494 1873 3497 1876 ne
rect 3497 1873 3552 1876
tri 3552 1873 3555 1876 sw
tri 3604 1873 3607 1876 ne
rect 3607 1873 3685 1876
tri 3685 1873 3689 1877 sw
tri 3497 1866 3504 1873 ne
rect 3504 1870 3555 1873
tri 3555 1870 3558 1873 sw
tri 3607 1870 3610 1873 ne
rect 3610 1870 3689 1873
rect 3504 1866 3558 1870
tri 3558 1866 3562 1870 sw
tri 3610 1866 3614 1870 ne
rect 3614 1866 3689 1870
tri 3689 1866 3696 1873 sw
rect 3236 1814 3242 1866
rect 3294 1814 3306 1866
rect 3358 1821 3434 1866
tri 3434 1821 3479 1866 sw
tri 3504 1821 3549 1866 ne
rect 3549 1821 3562 1866
tri 3562 1821 3607 1866 sw
tri 3614 1821 3659 1866 ne
rect 3659 1821 3696 1866
tri 3696 1821 3741 1866 sw
rect 3939 1821 3979 1906
rect 4887 1880 4893 1932
rect 4945 1880 4957 1932
rect 5009 1906 6572 1932
tri 6572 1906 6598 1932 sw
tri 6665 1906 6691 1932 ne
rect 6691 1906 11181 1932
tri 11181 1906 11219 1944 sw
rect 5009 1902 6598 1906
tri 6598 1902 6602 1906 sw
tri 6691 1902 6695 1906 ne
rect 6695 1902 11219 1906
rect 5009 1880 6602 1902
tri 6602 1880 6624 1902 sw
tri 11091 1880 11113 1902 ne
rect 11113 1880 11219 1902
tri 6550 1873 6557 1880 ne
rect 6557 1873 6624 1880
tri 6624 1873 6631 1880 sw
tri 11113 1873 11120 1880 ne
rect 11120 1873 11219 1880
tri 6557 1858 6572 1873 ne
rect 6572 1858 10594 1873
tri 6572 1843 6587 1858 ne
rect 6587 1843 10594 1858
tri 6587 1834 6596 1843 ne
rect 6596 1834 10594 1843
tri 3979 1821 3992 1834 sw
tri 6596 1833 6597 1834 ne
rect 6597 1833 10594 1834
rect 10588 1821 10594 1833
rect 10646 1821 10658 1873
rect 10710 1821 10716 1873
rect 10843 1821 10849 1873
rect 10901 1821 10913 1873
rect 10965 1871 11027 1873
tri 11027 1871 11029 1873 sw
tri 11120 1871 11122 1873 ne
rect 11122 1871 11219 1873
tri 11219 1871 11254 1906 sw
rect 10965 1845 11029 1871
tri 11029 1845 11055 1871 sw
tri 11122 1845 11148 1871 ne
rect 11148 1845 11254 1871
rect 10965 1843 11055 1845
tri 11055 1843 11057 1845 sw
tri 11148 1843 11150 1845 ne
rect 11150 1843 11254 1845
tri 11254 1843 11282 1871 sw
rect 13410 1859 13416 1871
tri 11896 1843 11912 1859 se
rect 11912 1843 13416 1859
rect 10965 1837 11057 1843
tri 11057 1837 11063 1843 sw
tri 11150 1837 11156 1843 ne
rect 11156 1837 11300 1843
rect 10965 1834 11063 1837
tri 11063 1834 11066 1837 sw
tri 11156 1834 11159 1837 ne
rect 11159 1834 11248 1837
rect 10965 1833 11066 1834
tri 11066 1833 11067 1834 sw
tri 11159 1833 11160 1834 ne
rect 11160 1833 11248 1834
rect 10965 1821 11067 1833
rect 3358 1814 3479 1821
tri 3479 1814 3486 1821 sw
tri 3549 1818 3552 1821 ne
rect 3552 1818 3607 1821
tri 3607 1818 3610 1821 sw
tri 3659 1818 3662 1821 ne
rect 3662 1818 3741 1821
tri 3552 1814 3556 1818 ne
rect 3556 1814 3610 1818
tri 3610 1814 3614 1818 sw
tri 3662 1814 3666 1818 ne
rect 3666 1814 3741 1818
tri 3741 1814 3748 1821 sw
rect 3939 1819 3992 1821
tri 3992 1819 3994 1821 sw
tri 11021 1819 11023 1821 ne
rect 11023 1819 11067 1821
tri 11067 1819 11081 1833 sw
tri 11160 1819 11174 1833 ne
rect 11174 1819 11248 1833
rect 3939 1816 3994 1819
tri 3939 1814 3941 1816 ne
rect 3941 1814 3994 1816
tri 3412 1792 3434 1814 ne
rect 3434 1793 3486 1814
tri 3486 1793 3507 1814 sw
tri 3556 1793 3577 1814 ne
rect 3577 1812 3614 1814
tri 3614 1812 3616 1814 sw
tri 3666 1812 3668 1814 ne
rect 3668 1812 3748 1814
rect 3577 1795 3616 1812
tri 3616 1795 3633 1812 sw
tri 3668 1795 3685 1812 ne
rect 3685 1795 3748 1812
tri 3748 1795 3767 1814 sw
tri 3941 1795 3960 1814 ne
rect 3960 1795 3994 1814
rect 3577 1793 3633 1795
tri 3633 1793 3635 1795 sw
tri 3685 1793 3687 1795 ne
rect 3687 1793 3767 1795
tri 3767 1793 3769 1795 sw
tri 3960 1793 3962 1795 ne
rect 3962 1793 3994 1795
tri 3994 1793 4020 1819 sw
tri 11023 1793 11049 1819 ne
rect 11049 1812 11081 1819
tri 11081 1812 11088 1819 sw
tri 11174 1812 11181 1819 ne
rect 11181 1812 11248 1819
rect 11049 1793 11088 1812
tri 11088 1793 11107 1812 sw
tri 11181 1793 11200 1812 ne
rect 11200 1793 11248 1812
rect 3434 1792 3507 1793
tri 3507 1792 3508 1793 sw
tri 3577 1792 3578 1793 ne
rect 3578 1792 3635 1793
tri 3635 1792 3636 1793 sw
tri 3687 1792 3688 1793 ne
rect 3688 1792 3769 1793
tri 3769 1792 3770 1793 sw
tri 3962 1792 3963 1793 ne
rect 3963 1792 10991 1793
tri 3434 1785 3441 1792 ne
rect 3441 1785 3508 1792
tri 3508 1785 3515 1792 sw
tri 3578 1785 3585 1792 ne
rect 3585 1785 3636 1792
tri 3636 1785 3643 1792 sw
tri 3688 1785 3695 1792 ne
rect 3695 1785 3770 1792
tri 3770 1785 3777 1792 sw
tri 3963 1785 3970 1792 ne
rect 3970 1786 10991 1792
tri 10991 1786 10998 1793 sw
tri 11049 1787 11055 1793 ne
rect 11055 1787 11107 1793
tri 11107 1787 11113 1793 sw
tri 11200 1787 11206 1793 ne
rect 11206 1787 11248 1793
tri 11055 1786 11056 1787 ne
rect 11056 1786 11113 1787
tri 11113 1786 11114 1787 sw
tri 11206 1786 11207 1787 ne
rect 11207 1786 11248 1787
rect 3970 1785 10998 1786
tri 10998 1785 10999 1786 sw
tri 11056 1785 11057 1786 ne
rect 11057 1785 11114 1786
tri 11114 1785 11115 1786 sw
tri 11207 1785 11208 1786 ne
rect 11208 1785 11248 1786
tri 11872 1819 11896 1843 se
rect 11896 1819 13416 1843
rect 13468 1819 13480 1871
rect 13532 1819 13538 1871
tri 11854 1801 11872 1819 se
rect 11872 1801 11912 1819
tri 11912 1801 11930 1819 nw
tri 11839 1786 11854 1801 se
rect 11854 1786 11897 1801
tri 11897 1786 11912 1801 nw
tri 3441 1773 3453 1785 ne
rect 3453 1776 3515 1785
tri 3515 1776 3524 1785 sw
tri 3585 1776 3594 1785 ne
rect 3594 1776 3643 1785
tri 3643 1776 3652 1785 sw
tri 3695 1776 3704 1785 ne
rect 3704 1776 3777 1785
tri 3777 1776 3786 1785 sw
tri 3970 1776 3979 1785 ne
rect 3979 1776 10999 1785
rect 3453 1773 3524 1776
tri 3524 1773 3527 1776 sw
tri 3594 1773 3597 1776 ne
rect 3597 1773 3652 1776
tri 3652 1773 3655 1776 sw
tri 3704 1773 3707 1776 ne
rect 3707 1773 3786 1776
tri 3786 1773 3789 1776 sw
tri 3979 1773 3982 1776 ne
rect 3982 1773 10999 1776
tri 10999 1773 11011 1785 sw
tri 11057 1773 11069 1785 ne
rect 11069 1781 11115 1785
tri 11115 1781 11119 1785 sw
tri 11208 1781 11212 1785 ne
rect 11212 1781 11300 1785
rect 11069 1773 11119 1781
tri 11119 1773 11127 1781 sw
rect 11248 1773 11300 1781
tri 3453 1721 3505 1773 ne
rect 3505 1765 3527 1773
tri 3527 1765 3535 1773 sw
tri 3597 1765 3605 1773 ne
rect 3605 1765 3655 1773
tri 3655 1765 3663 1773 sw
tri 3707 1765 3715 1773 ne
rect 3715 1765 3789 1773
tri 3789 1765 3797 1773 sw
tri 3982 1765 3990 1773 ne
rect 3990 1765 11011 1773
tri 11011 1765 11019 1773 sw
tri 11069 1765 11077 1773 ne
rect 11077 1765 11127 1773
tri 11127 1765 11135 1773 sw
rect 3505 1753 3535 1765
tri 3535 1753 3547 1765 sw
tri 3605 1760 3610 1765 ne
rect 3610 1760 3663 1765
tri 3663 1760 3668 1765 sw
tri 3715 1760 3720 1765 ne
rect 3720 1760 3797 1765
tri 3610 1753 3617 1760 ne
rect 3617 1754 3668 1760
tri 3668 1754 3674 1760 sw
tri 3720 1754 3726 1760 ne
rect 3726 1754 3797 1760
rect 3617 1753 3674 1754
tri 3674 1753 3675 1754 sw
tri 3726 1753 3727 1754 ne
rect 3727 1753 3797 1754
tri 3797 1753 3809 1765 sw
tri 3990 1753 4002 1765 ne
rect 4002 1753 11019 1765
rect 3505 1721 3547 1753
tri 3547 1721 3579 1753 sw
tri 3617 1721 3649 1753 ne
rect 3649 1721 3675 1753
tri 3675 1721 3707 1753 sw
tri 3727 1721 3759 1753 ne
rect 3759 1721 3809 1753
tri 3809 1721 3841 1753 sw
tri 10973 1721 11005 1753 ne
rect 11005 1729 11019 1753
tri 11019 1729 11055 1765 sw
tri 11077 1729 11113 1765 ne
rect 11113 1729 11135 1765
tri 11135 1729 11171 1765 sw
rect 11005 1728 11055 1729
tri 11055 1728 11056 1729 sw
tri 11113 1728 11114 1729 ne
rect 11114 1728 11171 1729
tri 11171 1728 11172 1729 sw
rect 11005 1721 11056 1728
tri 11056 1721 11063 1728 sw
tri 11114 1721 11121 1728 ne
rect 11121 1721 11172 1728
tri 11172 1721 11179 1728 sw
tri 11796 1743 11839 1786 se
rect 11839 1743 11854 1786
tri 11854 1743 11897 1786 nw
tri 11912 1743 11955 1786 se
rect 11955 1746 13473 1786
rect 11955 1743 11961 1746
tri 11787 1734 11796 1743 se
rect 11796 1734 11845 1743
tri 11845 1734 11854 1743 nw
tri 11903 1734 11912 1743 se
rect 11912 1734 11961 1743
tri 11961 1734 11973 1746 nw
rect 13467 1734 13473 1746
rect 13525 1734 13537 1786
rect 13589 1734 13595 1786
tri 11781 1728 11787 1734 se
rect 11787 1728 11839 1734
tri 11839 1728 11845 1734 nw
tri 11897 1728 11903 1734 se
rect 11903 1728 11955 1734
tri 11955 1728 11961 1734 nw
tri 3505 1720 3506 1721 ne
rect 3506 1720 3579 1721
tri 3579 1720 3580 1721 sw
tri 3649 1720 3650 1721 ne
rect 3650 1720 3707 1721
tri 3707 1720 3708 1721 sw
tri 3759 1720 3760 1721 ne
rect 3760 1720 3841 1721
tri 3841 1720 3842 1721 sw
tri 11005 1720 11006 1721 ne
rect 11006 1720 11063 1721
tri 3506 1718 3508 1720 ne
rect 3508 1718 3580 1720
tri 3580 1718 3582 1720 sw
tri 3650 1718 3652 1720 ne
rect 3652 1718 3708 1720
tri 3708 1718 3710 1720 sw
tri 3760 1718 3762 1720 ne
rect 3762 1718 3842 1720
tri 3842 1718 3844 1720 sw
tri 3508 1668 3558 1718 ne
rect 3558 1713 3582 1718
tri 3582 1713 3587 1718 sw
tri 3652 1713 3657 1718 ne
rect 3657 1713 3710 1718
tri 3710 1713 3715 1718 sw
tri 3762 1713 3767 1718 ne
rect 3767 1713 3844 1718
tri 3844 1713 3849 1718 sw
rect 3558 1702 3587 1713
tri 3587 1702 3598 1713 sw
tri 3657 1702 3668 1713 ne
rect 3668 1702 3715 1713
tri 3715 1702 3726 1713 sw
tri 3767 1702 3778 1713 ne
rect 3778 1702 10482 1713
rect 3558 1673 3598 1702
tri 3598 1673 3627 1702 sw
tri 3668 1673 3697 1702 ne
rect 3697 1696 3726 1702
tri 3726 1696 3732 1702 sw
tri 3778 1696 3784 1702 ne
rect 3784 1696 10482 1702
rect 3697 1673 3732 1696
tri 3732 1673 3755 1696 sw
tri 3784 1673 3807 1696 ne
rect 3807 1673 10482 1696
tri 10482 1673 10522 1713 sw
rect 3558 1668 3627 1673
tri 3627 1668 3632 1673 sw
tri 3697 1668 3702 1673 ne
rect 3702 1668 3755 1673
tri 3755 1668 3760 1673 sw
tri 10448 1668 10453 1673 ne
rect 10453 1668 10522 1673
tri 10522 1668 10527 1673 sw
rect 10578 1668 10584 1720
rect 10636 1668 10648 1720
rect 10700 1713 10706 1720
tri 11006 1713 11013 1720 ne
rect 11013 1713 11063 1720
rect 10700 1707 10969 1713
tri 10969 1707 10975 1713 sw
tri 11013 1707 11019 1713 ne
rect 11019 1707 11063 1713
tri 11063 1707 11077 1721 sw
tri 11121 1707 11135 1721 ne
rect 11135 1715 11179 1721
tri 11179 1715 11185 1721 sw
rect 11248 1715 11300 1721
tri 11768 1715 11781 1728 se
rect 11781 1715 11817 1728
rect 11135 1707 11185 1715
tri 11185 1707 11193 1715 sw
tri 11760 1707 11768 1715 se
rect 11768 1707 11817 1715
rect 10700 1706 10975 1707
tri 10975 1706 10976 1707 sw
tri 11019 1706 11020 1707 ne
rect 11020 1706 11077 1707
tri 11077 1706 11078 1707 sw
tri 11135 1706 11136 1707 ne
rect 11136 1706 11193 1707
tri 11193 1706 11194 1707 sw
tri 11759 1706 11760 1707 se
rect 11760 1706 11817 1707
tri 11817 1706 11839 1728 nw
tri 11875 1706 11897 1728 se
rect 11897 1706 11933 1728
tri 11933 1706 11955 1728 nw
rect 10700 1680 10976 1706
tri 10976 1680 11002 1706 sw
tri 11020 1680 11046 1706 ne
rect 11046 1680 11078 1706
rect 10700 1673 11002 1680
rect 10700 1668 10706 1673
tri 10952 1668 10957 1673 ne
rect 10957 1668 11002 1673
tri 3558 1654 3572 1668 ne
rect 3572 1654 3632 1668
tri 3632 1654 3646 1668 sw
tri 3702 1654 3716 1668 ne
rect 3716 1654 3760 1668
tri 3760 1654 3774 1668 sw
tri 10453 1654 10467 1668 ne
rect 10467 1654 10527 1668
tri 10527 1654 10541 1668 sw
tri 10957 1654 10971 1668 ne
rect 10971 1667 11002 1668
tri 11002 1667 11015 1680 sw
tri 11046 1667 11059 1680 ne
rect 11059 1671 11078 1680
tri 11078 1671 11113 1706 sw
tri 11136 1671 11171 1706 ne
rect 11171 1685 11194 1706
tri 11194 1685 11215 1706 sw
tri 11738 1685 11759 1706 se
rect 11759 1685 11796 1706
tri 11796 1685 11817 1706 nw
tri 11854 1685 11875 1706 se
rect 11875 1685 11897 1706
rect 11171 1671 11215 1685
tri 11215 1671 11229 1685 sw
tri 11724 1671 11738 1685 se
rect 11738 1671 11781 1685
rect 11059 1670 11113 1671
tri 11113 1670 11114 1671 sw
tri 11171 1670 11172 1671 ne
rect 11172 1670 11229 1671
tri 11229 1670 11230 1671 sw
tri 11723 1670 11724 1671 se
rect 11724 1670 11781 1671
tri 11781 1670 11796 1685 nw
tri 11839 1670 11854 1685 se
rect 11854 1670 11897 1685
tri 11897 1670 11933 1706 nw
tri 11955 1670 11991 1706 se
rect 11991 1670 13473 1706
rect 11059 1667 11114 1670
rect 10971 1654 11015 1667
tri 11015 1654 11028 1667 sw
tri 11059 1654 11072 1667 ne
rect 11072 1654 11114 1667
tri 11114 1654 11130 1670 sw
tri 11172 1654 11188 1670 ne
rect 11188 1654 11230 1670
tri 11230 1654 11246 1670 sw
tri 11707 1654 11723 1670 se
rect 11723 1654 11765 1670
tri 11765 1654 11781 1670 nw
tri 11823 1654 11839 1670 se
rect 11839 1654 11881 1670
tri 11881 1654 11897 1670 nw
tri 11939 1654 11955 1670 se
rect 11955 1666 13473 1670
rect 11955 1654 11997 1666
tri 11997 1654 12009 1666 nw
tri 13316 1654 13328 1666 ne
rect 13328 1654 13473 1666
rect 13525 1654 13537 1706
rect 13589 1654 13595 1706
tri 3572 1649 3577 1654 ne
rect 3577 1649 3646 1654
rect 2767 1593 2776 1649
rect 2832 1593 2859 1649
rect 2915 1630 2941 1649
rect 2997 1630 3006 1649
tri 3577 1644 3582 1649 ne
rect 3582 1644 3646 1649
tri 3646 1644 3656 1654 sw
tri 3716 1644 3726 1654 ne
rect 3726 1644 3774 1654
tri 3774 1644 3784 1654 sw
tri 10467 1644 10477 1654 ne
rect 10477 1644 10541 1654
tri 3582 1643 3583 1644 ne
rect 3583 1643 3656 1644
tri 3656 1643 3657 1644 sw
tri 3726 1643 3727 1644 ne
rect 3727 1643 6346 1644
tri 6346 1643 6347 1644 sw
tri 10477 1643 10478 1644 ne
rect 10478 1643 10541 1644
tri 3583 1630 3596 1643 ne
rect 3596 1630 3657 1643
rect 2916 1593 2941 1630
rect 2767 1578 2779 1593
rect 2831 1578 2864 1593
rect 2916 1578 2949 1593
rect 3001 1578 3007 1630
tri 3596 1591 3635 1630 ne
rect 3635 1591 3657 1630
tri 3657 1591 3709 1643 sw
tri 3727 1635 3735 1643 ne
rect 3735 1635 6347 1643
tri 6347 1635 6355 1643 sw
tri 3735 1602 3768 1635 ne
rect 3768 1602 6355 1635
tri 6330 1591 6341 1602 ne
rect 6341 1591 6355 1602
tri 6355 1591 6399 1635 sw
rect 7685 1591 7691 1643
rect 7743 1591 7755 1643
rect 7807 1633 7813 1643
tri 10478 1639 10482 1643 ne
rect 10482 1639 10541 1643
tri 10541 1639 10556 1654 sw
tri 10971 1639 10986 1654 ne
rect 10986 1649 11028 1654
tri 11028 1649 11033 1654 sw
tri 11072 1649 11077 1654 ne
rect 11077 1649 11130 1654
tri 11130 1649 11135 1654 sw
tri 11188 1649 11193 1654 ne
rect 11193 1649 11246 1654
tri 11246 1649 11251 1654 sw
tri 11702 1649 11707 1654 se
rect 11707 1649 11738 1654
rect 10986 1639 11033 1649
tri 10482 1633 10488 1639 ne
rect 10488 1633 10820 1639
rect 7807 1598 10356 1633
tri 10356 1598 10391 1633 sw
tri 10488 1623 10498 1633 ne
rect 10498 1623 10820 1633
tri 10498 1598 10523 1623 ne
rect 10523 1598 10820 1623
rect 7807 1593 10391 1598
rect 7807 1591 7813 1593
tri 10338 1591 10340 1593 ne
rect 10340 1591 10391 1593
tri 10391 1591 10398 1598 sw
tri 10523 1591 10530 1598 ne
rect 10530 1591 10820 1598
tri 3635 1587 3639 1591 ne
rect 3639 1587 3709 1591
tri 3709 1587 3713 1591 sw
tri 6341 1587 6345 1591 ne
rect 6345 1587 6399 1591
tri 6399 1587 6403 1591 sw
tri 10340 1587 10344 1591 ne
rect 10344 1587 10398 1591
tri 10398 1587 10402 1591 sw
tri 10530 1587 10534 1591 ne
rect 10534 1587 10820 1591
rect 10872 1587 10884 1639
rect 10936 1587 10942 1639
tri 10986 1633 10992 1639 ne
rect 10992 1633 11033 1639
tri 11033 1633 11049 1649 sw
tri 11077 1633 11093 1649 ne
rect 11093 1633 11135 1649
tri 10992 1626 10999 1633 ne
rect 10999 1626 11049 1633
tri 11049 1626 11056 1633 sw
tri 11093 1626 11100 1633 ne
rect 11100 1626 11135 1633
tri 11135 1626 11158 1649 sw
tri 11193 1626 11216 1649 ne
rect 11216 1627 11251 1649
tri 11251 1627 11273 1649 sw
tri 11680 1627 11702 1649 se
rect 11702 1627 11738 1649
tri 11738 1627 11765 1654 nw
tri 11796 1627 11823 1654 se
rect 11823 1648 11875 1654
tri 11875 1648 11881 1654 nw
tri 11933 1648 11939 1654 se
rect 11939 1648 11991 1654
tri 11991 1648 11997 1654 nw
rect 11823 1627 11853 1648
rect 11216 1626 11273 1627
tri 11273 1626 11274 1627 sw
tri 11679 1626 11680 1627 se
rect 11680 1626 11737 1627
tri 11737 1626 11738 1627 nw
tri 11795 1626 11796 1627 se
rect 11796 1626 11853 1627
tri 11853 1626 11875 1648 nw
tri 11911 1626 11933 1648 se
rect 11933 1626 11969 1648
tri 11969 1626 11991 1648 nw
tri 10999 1623 11002 1626 ne
rect 11002 1623 11056 1626
tri 11056 1623 11059 1626 sw
tri 11100 1623 11103 1626 ne
rect 11103 1623 11158 1626
tri 11002 1598 11027 1623 ne
rect 11027 1610 11059 1623
tri 11059 1610 11072 1623 sw
tri 11103 1610 11116 1623 ne
rect 11116 1613 11158 1623
tri 11158 1613 11171 1626 sw
tri 11216 1613 11229 1626 ne
rect 11229 1613 11274 1626
tri 11274 1613 11287 1626 sw
tri 11666 1613 11679 1626 se
rect 11679 1613 11723 1626
rect 11116 1612 11171 1613
tri 11171 1612 11172 1613 sw
tri 11229 1612 11230 1613 ne
rect 11230 1612 11287 1613
tri 11287 1612 11288 1613 sw
tri 11665 1612 11666 1613 se
rect 11666 1612 11723 1613
tri 11723 1612 11737 1626 nw
tri 11781 1612 11795 1626 se
rect 11795 1612 11839 1626
tri 11839 1612 11853 1626 nw
tri 11897 1612 11911 1626 se
rect 11911 1612 11955 1626
tri 11955 1612 11969 1626 nw
tri 12013 1612 12027 1626 se
rect 12027 1612 14225 1626
rect 11116 1610 11172 1612
rect 11027 1598 11072 1610
tri 11072 1598 11084 1610 sw
tri 11116 1598 11128 1610 ne
rect 11128 1598 11172 1610
tri 11027 1591 11034 1598 ne
rect 11034 1591 11084 1598
tri 11084 1591 11091 1598 sw
tri 11128 1591 11135 1598 ne
rect 11135 1591 11172 1598
tri 11172 1591 11193 1612 sw
tri 11230 1591 11251 1612 ne
rect 11251 1591 11288 1612
tri 11288 1591 11309 1612 sw
tri 11644 1591 11665 1612 se
rect 11665 1591 11685 1612
tri 11034 1587 11038 1591 ne
rect 11038 1587 11091 1591
rect 2767 1559 3007 1578
tri 3639 1574 3652 1587 ne
rect 3652 1574 3713 1587
tri 3713 1574 3726 1587 sw
tri 6345 1577 6355 1587 ne
rect 6355 1577 6403 1587
tri 6403 1577 6413 1587 sw
tri 10344 1577 10354 1587 ne
rect 10354 1577 10402 1587
tri 6355 1574 6358 1577 ne
rect 6358 1574 6413 1577
tri 6413 1574 6416 1577 sw
tri 10354 1574 10357 1577 ne
rect 10357 1574 10402 1577
tri 10402 1574 10415 1587 sw
tri 11038 1574 11051 1587 ne
rect 11051 1574 11091 1587
tri 11091 1574 11108 1591 sw
tri 11135 1574 11152 1591 ne
rect 11152 1574 11193 1591
tri 11193 1574 11210 1591 sw
tri 11251 1574 11268 1591 ne
rect 11268 1574 11309 1591
tri 11309 1574 11326 1591 sw
tri 11627 1574 11644 1591 se
rect 11644 1574 11685 1591
tri 11685 1574 11723 1612 nw
tri 11743 1574 11781 1612 se
rect 11781 1590 11817 1612
tri 11817 1590 11839 1612 nw
tri 11875 1590 11897 1612 se
rect 11897 1590 11933 1612
tri 11933 1590 11955 1612 nw
tri 11991 1590 12013 1612 se
rect 12013 1590 14225 1612
rect 11781 1574 11801 1590
tri 11801 1574 11817 1590 nw
tri 11859 1574 11875 1590 se
rect 11875 1574 11917 1590
tri 11917 1574 11933 1590 nw
tri 11975 1574 11991 1590 se
rect 11991 1586 14225 1590
rect 11991 1574 12033 1586
tri 12033 1574 12045 1586 nw
rect 14219 1574 14225 1586
rect 14277 1574 14289 1626
rect 14341 1574 14347 1626
tri 3652 1570 3656 1574 ne
rect 3656 1570 3726 1574
tri 3726 1570 3730 1574 sw
tri 6358 1570 6362 1574 ne
rect 6362 1570 6416 1574
tri 6416 1570 6420 1574 sw
tri 10357 1570 10361 1574 ne
rect 10361 1570 10415 1574
rect 2767 1503 2776 1559
rect 2832 1503 2859 1559
rect 2915 1558 2941 1559
rect 2997 1558 3007 1559
rect 2916 1506 2941 1558
rect 3001 1506 3007 1558
tri 3656 1552 3674 1570 ne
rect 3674 1552 3730 1570
tri 3730 1552 3748 1570 sw
tri 6362 1552 6380 1570 ne
rect 6380 1552 6420 1570
tri 6420 1552 6438 1570 sw
tri 10361 1552 10379 1570 ne
rect 10379 1552 10415 1570
tri 3674 1540 3686 1552 ne
rect 3686 1540 4455 1552
tri 3686 1506 3720 1540 ne
rect 3720 1506 4455 1540
rect 2915 1503 2941 1506
rect 2997 1503 3006 1506
tri 3720 1503 3723 1506 ne
rect 3723 1503 4455 1506
tri 3723 1500 3726 1503 ne
rect 3726 1500 4455 1503
rect 4507 1500 4525 1552
rect 4577 1500 4595 1552
rect 4647 1500 4665 1552
rect 4717 1500 4735 1552
rect 4787 1500 4805 1552
rect 4857 1500 4875 1552
rect 4927 1500 4944 1552
rect 4996 1500 5002 1552
tri 6380 1519 6413 1552 ne
rect 6413 1540 6438 1552
tri 6438 1540 6450 1552 sw
tri 10379 1540 10391 1552 ne
rect 10391 1540 10415 1552
tri 10415 1540 10449 1574 sw
tri 11051 1566 11059 1574 ne
rect 11059 1566 11108 1574
tri 11108 1566 11116 1574 sw
tri 11152 1566 11160 1574 ne
rect 11160 1566 11210 1574
tri 11059 1540 11085 1566 ne
rect 11085 1553 11116 1566
tri 11116 1553 11129 1566 sw
tri 11160 1553 11173 1566 ne
rect 11173 1555 11210 1566
tri 11210 1555 11229 1574 sw
tri 11268 1555 11287 1574 ne
rect 11287 1569 11326 1574
tri 11326 1569 11331 1574 sw
tri 11622 1569 11627 1574 se
rect 11627 1569 11680 1574
tri 11680 1569 11685 1574 nw
tri 11738 1569 11743 1574 se
rect 11743 1569 11781 1574
rect 11287 1555 11331 1569
tri 11331 1555 11345 1569 sw
tri 11608 1555 11622 1569 se
rect 11622 1555 11666 1569
tri 11666 1555 11680 1569 nw
tri 11724 1555 11738 1569 se
rect 11738 1555 11781 1569
rect 11173 1554 11229 1555
tri 11229 1554 11230 1555 sw
tri 11287 1554 11288 1555 ne
rect 11288 1554 11665 1555
tri 11665 1554 11666 1555 nw
tri 11723 1554 11724 1555 se
rect 11724 1554 11781 1555
tri 11781 1554 11801 1574 nw
tri 11853 1568 11859 1574 se
rect 11859 1568 11911 1574
tri 11911 1568 11917 1574 nw
tri 11969 1568 11975 1574 se
rect 11975 1568 12027 1574
tri 12027 1568 12033 1574 nw
tri 11839 1554 11853 1568 se
rect 11853 1554 11897 1568
tri 11897 1554 11911 1568 nw
tri 11955 1554 11969 1568 se
rect 11173 1553 11230 1554
rect 11085 1540 11129 1553
tri 11129 1540 11142 1553 sw
tri 11173 1540 11186 1553 ne
rect 11186 1540 11230 1553
rect 6413 1519 6450 1540
tri 6450 1519 6471 1540 sw
tri 10391 1519 10412 1540 ne
rect 10412 1533 11012 1540
tri 11012 1533 11019 1540 sw
tri 11085 1533 11092 1540 ne
rect 11092 1533 11142 1540
tri 11142 1533 11149 1540 sw
tri 11186 1533 11193 1540 ne
rect 11193 1533 11230 1540
tri 11230 1533 11251 1554 sw
tri 11288 1533 11309 1554 ne
rect 11309 1533 11626 1554
rect 10412 1519 11019 1533
tri 6413 1500 6432 1519 ne
rect 6432 1500 6471 1519
tri 6471 1500 6490 1519 sw
tri 10412 1500 10431 1519 ne
rect 10431 1509 11019 1519
tri 11019 1509 11043 1533 sw
tri 11092 1509 11116 1533 ne
rect 11116 1509 11149 1533
tri 11149 1509 11173 1533 sw
tri 11193 1509 11217 1533 ne
rect 11217 1515 11251 1533
tri 11251 1515 11269 1533 sw
tri 11309 1515 11327 1533 ne
rect 11327 1515 11626 1533
tri 11626 1515 11665 1554 nw
tri 11684 1515 11723 1554 se
rect 11723 1532 11759 1554
tri 11759 1532 11781 1554 nw
tri 11817 1532 11839 1554 se
rect 11839 1532 11875 1554
tri 11875 1532 11897 1554 nw
tri 11933 1532 11955 1554 se
rect 11955 1532 11969 1554
rect 11217 1509 11269 1515
rect 10431 1500 11043 1509
tri 6432 1461 6471 1500 ne
rect 6471 1489 6490 1500
tri 6490 1489 6501 1500 sw
tri 10994 1489 11005 1500 ne
rect 11005 1489 11043 1500
tri 11043 1489 11063 1509 sw
tri 11116 1489 11136 1509 ne
rect 11136 1496 11173 1509
tri 11173 1496 11186 1509 sw
tri 11217 1496 11230 1509 ne
rect 11230 1496 11269 1509
tri 11269 1496 11288 1515 sw
tri 11665 1496 11684 1515 se
rect 11684 1496 11723 1515
tri 11723 1496 11759 1532 nw
tri 11795 1510 11817 1532 se
rect 11817 1510 11853 1532
tri 11853 1510 11875 1532 nw
tri 11911 1510 11933 1532 se
rect 11933 1510 11969 1532
tri 11969 1510 12027 1568 nw
tri 11781 1496 11795 1510 se
rect 11795 1496 11839 1510
tri 11839 1496 11853 1510 nw
tri 11897 1496 11911 1510 se
rect 11136 1489 11186 1496
tri 11186 1489 11193 1496 sw
tri 11230 1489 11237 1496 ne
rect 11237 1489 11288 1496
rect 6471 1482 6501 1489
tri 6501 1482 6508 1489 sw
tri 11005 1482 11012 1489 ne
rect 11012 1482 11063 1489
rect 6471 1461 6508 1482
tri 6508 1461 6529 1482 sw
tri 11012 1461 11033 1482 ne
rect 11033 1475 11063 1482
tri 11063 1475 11077 1489 sw
tri 11136 1475 11150 1489 ne
rect 11150 1475 11193 1489
tri 11193 1475 11207 1489 sw
tri 11237 1475 11251 1489 ne
rect 11251 1475 11288 1489
tri 11288 1475 11309 1496 sw
tri 11644 1475 11665 1496 se
rect 11665 1475 11702 1496
tri 11702 1475 11723 1496 nw
tri 11760 1475 11781 1496 se
rect 11781 1475 11818 1496
tri 11818 1475 11839 1496 nw
tri 11876 1475 11897 1496 se
rect 11897 1475 11911 1496
rect 11033 1461 11077 1475
tri 6471 1452 6480 1461 ne
rect 6480 1458 10706 1461
tri 10706 1458 10709 1461 sw
tri 11033 1458 11036 1461 ne
rect 11036 1458 11077 1461
rect 6480 1452 10709 1458
tri 10709 1452 10715 1458 sw
rect 10820 1452 10872 1458
tri 6480 1447 6485 1452 ne
rect 6485 1447 10715 1452
tri 10715 1447 10720 1452 sw
tri 6485 1419 6513 1447 ne
rect 6513 1419 10820 1447
tri 10690 1400 10709 1419 ne
rect 10709 1400 10820 1419
tri 11036 1431 11063 1458 ne
rect 11063 1452 11077 1458
tri 11077 1452 11100 1475 sw
tri 11150 1452 11173 1475 ne
rect 11173 1452 11207 1475
tri 11207 1452 11230 1475 sw
tri 11251 1452 11274 1475 ne
rect 11274 1474 11701 1475
tri 11701 1474 11702 1475 nw
tri 11759 1474 11760 1475 se
rect 11760 1474 11817 1475
tri 11817 1474 11818 1475 nw
tri 11875 1474 11876 1475 se
rect 11876 1474 11911 1475
rect 11274 1452 11662 1474
rect 11063 1435 11100 1452
tri 11100 1435 11117 1452 sw
tri 11173 1435 11190 1452 ne
rect 11190 1439 11230 1452
tri 11230 1439 11243 1452 sw
tri 11274 1439 11287 1452 ne
rect 11287 1439 11662 1452
rect 11190 1435 11243 1439
tri 11243 1435 11247 1439 sw
tri 11287 1435 11291 1439 ne
rect 11291 1435 11662 1439
tri 11662 1435 11701 1474 nw
tri 11737 1452 11759 1474 se
rect 11759 1452 11795 1474
tri 11795 1452 11817 1474 nw
tri 11853 1452 11875 1474 se
rect 11875 1452 11911 1474
tri 11911 1452 11969 1510 nw
tri 11720 1435 11737 1452 se
rect 11737 1435 11778 1452
tri 11778 1435 11795 1452 nw
tri 11836 1435 11853 1452 se
rect 11063 1431 11117 1435
tri 11117 1431 11121 1435 sw
tri 11190 1431 11194 1435 ne
rect 11194 1431 11247 1435
tri 11247 1431 11251 1435 sw
tri 11716 1431 11720 1435 se
rect 11720 1431 11759 1435
rect 10820 1388 10872 1400
tri 11063 1373 11121 1431 ne
tri 11121 1394 11158 1431 sw
tri 11194 1395 11230 1431 ne
rect 11230 1416 11251 1431
tri 11251 1416 11266 1431 sw
tri 11701 1416 11716 1431 se
rect 11716 1416 11759 1431
tri 11759 1416 11778 1435 nw
tri 11817 1416 11836 1435 se
rect 11836 1416 11853 1435
rect 11230 1395 11266 1416
tri 11266 1395 11287 1416 sw
tri 11680 1395 11701 1416 se
rect 11701 1395 11738 1416
tri 11738 1395 11759 1416 nw
tri 11796 1395 11817 1416 se
rect 11817 1395 11853 1416
tri 11230 1394 11231 1395 ne
rect 11231 1394 11737 1395
tri 11737 1394 11738 1395 nw
tri 11795 1394 11796 1395 se
rect 11796 1394 11853 1395
tri 11853 1394 11911 1452 nw
rect 11121 1373 11158 1394
tri 11158 1373 11179 1394 sw
tri 11231 1373 11252 1394 ne
rect 11252 1373 11698 1394
rect 10820 1330 10872 1336
tri 11121 1330 11164 1373 ne
rect 11164 1336 11179 1373
tri 11179 1336 11216 1373 sw
tri 11252 1355 11270 1373 ne
rect 11270 1355 11698 1373
tri 11698 1355 11737 1394 nw
tri 11756 1355 11795 1394 se
tri 11737 1336 11756 1355 se
rect 11756 1336 11795 1355
tri 11795 1336 11853 1394 nw
rect 11164 1330 11216 1336
tri 11164 1315 11179 1330 ne
rect 11179 1315 11216 1330
tri 11216 1315 11237 1336 sw
tri 11716 1315 11737 1336 se
rect 11737 1315 11774 1336
tri 11774 1315 11795 1336 nw
tri 11179 1275 11219 1315 ne
rect 11219 1275 11734 1315
tri 11734 1275 11774 1315 nw
<< via2 >>
rect 2788 2731 2844 2732
rect 2874 2731 2930 2732
rect 2960 2731 3016 2732
rect 3046 2731 3102 2732
rect 3131 2731 3187 2732
rect 3216 2731 3272 2732
rect 3301 2731 3357 2732
rect 3386 2731 3442 2732
rect 2788 2679 2793 2731
rect 2793 2679 2844 2731
rect 2874 2679 2892 2731
rect 2892 2679 2930 2731
rect 2960 2679 2991 2731
rect 2991 2679 3016 2731
rect 3046 2679 3089 2731
rect 3089 2679 3102 2731
rect 3131 2679 3141 2731
rect 3141 2679 3187 2731
rect 3216 2679 3239 2731
rect 3239 2679 3272 2731
rect 3301 2679 3337 2731
rect 3337 2679 3357 2731
rect 3386 2679 3435 2731
rect 3435 2679 3442 2731
rect 2788 2676 2844 2679
rect 2874 2676 2930 2679
rect 2960 2676 3016 2679
rect 3046 2676 3102 2679
rect 3131 2676 3187 2679
rect 3216 2676 3272 2679
rect 3301 2676 3357 2679
rect 3386 2676 3442 2679
rect 3471 2731 3527 2732
rect 3471 2679 3481 2731
rect 3481 2679 3527 2731
rect 3471 2676 3527 2679
rect 2788 2643 2844 2648
rect 2874 2643 2930 2648
rect 2960 2643 3016 2648
rect 3046 2643 3102 2648
rect 3131 2643 3187 2648
rect 3216 2643 3272 2648
rect 3301 2643 3357 2648
rect 3386 2643 3442 2648
rect 2788 2592 2793 2643
rect 2793 2592 2844 2643
rect 2874 2592 2892 2643
rect 2892 2592 2930 2643
rect 2960 2592 2991 2643
rect 2991 2592 3016 2643
rect 3046 2592 3089 2643
rect 3089 2592 3102 2643
rect 3131 2592 3141 2643
rect 3141 2592 3187 2643
rect 3216 2592 3239 2643
rect 3239 2592 3272 2643
rect 3301 2592 3337 2643
rect 3337 2592 3357 2643
rect 3386 2592 3435 2643
rect 3435 2592 3442 2643
rect 3471 2643 3527 2648
rect 3471 2592 3481 2643
rect 3481 2592 3527 2643
rect 2788 2555 2844 2564
rect 2874 2555 2930 2564
rect 2960 2555 3016 2564
rect 3046 2555 3102 2564
rect 3131 2555 3187 2564
rect 3216 2555 3272 2564
rect 3301 2555 3357 2564
rect 3386 2555 3442 2564
rect 2788 2508 2793 2555
rect 2793 2508 2844 2555
rect 2874 2508 2892 2555
rect 2892 2508 2930 2555
rect 2960 2508 2991 2555
rect 2991 2508 3016 2555
rect 3046 2508 3089 2555
rect 3089 2508 3102 2555
rect 3131 2508 3141 2555
rect 3141 2508 3187 2555
rect 3216 2508 3239 2555
rect 3239 2508 3272 2555
rect 3301 2508 3337 2555
rect 3337 2508 3357 2555
rect 3386 2508 3435 2555
rect 3435 2508 3442 2555
rect 3471 2555 3527 2564
rect 3471 2508 3481 2555
rect 3481 2508 3527 2555
rect 2776 1630 2832 1649
rect 2776 1593 2779 1630
rect 2779 1593 2831 1630
rect 2831 1593 2832 1630
rect 2859 1630 2915 1649
rect 2941 1630 2997 1649
rect 2859 1593 2864 1630
rect 2864 1593 2915 1630
rect 2941 1593 2949 1630
rect 2949 1593 2997 1630
rect 2776 1558 2832 1559
rect 2776 1506 2779 1558
rect 2779 1506 2831 1558
rect 2831 1506 2832 1558
rect 2776 1503 2832 1506
rect 2859 1558 2915 1559
rect 2941 1558 2997 1559
rect 2859 1506 2864 1558
rect 2864 1506 2915 1558
rect 2941 1506 2949 1558
rect 2949 1506 2997 1558
rect 2859 1503 2915 1506
rect 2941 1503 2997 1506
<< metal3 >>
tri 2771 2761 3000 2990 se
rect 3000 2761 3545 2895
rect 2771 2732 3545 2761
rect 2771 2676 2788 2732
rect 2844 2676 2874 2732
rect 2930 2676 2960 2732
rect 3016 2676 3046 2732
rect 3102 2676 3131 2732
rect 3187 2676 3216 2732
rect 3272 2676 3301 2732
rect 3357 2676 3386 2732
rect 3442 2676 3471 2732
rect 3527 2676 3545 2732
rect 2771 2648 3545 2676
rect 2771 2592 2788 2648
rect 2844 2592 2874 2648
rect 2930 2592 2960 2648
rect 3016 2592 3046 2648
rect 3102 2592 3131 2648
rect 3187 2592 3216 2648
rect 3272 2592 3301 2648
rect 3357 2592 3386 2648
rect 3442 2592 3471 2648
rect 3527 2592 3545 2648
rect 2771 2564 3545 2592
rect 2771 2508 2788 2564
rect 2844 2508 2874 2564
rect 2930 2508 2960 2564
rect 3016 2508 3046 2564
rect 3102 2508 3131 2564
rect 3187 2508 3216 2564
rect 3272 2508 3301 2564
rect 3357 2508 3386 2564
rect 3442 2508 3471 2564
rect 3527 2508 3545 2564
rect 2771 2497 3545 2508
rect 2771 1649 3009 2497
tri 3009 2400 3106 2497 nw
rect 2771 1593 2776 1649
rect 2832 1593 2859 1649
rect 2915 1593 2941 1649
rect 2997 1593 3009 1649
rect 2771 1559 3009 1593
rect 2771 1503 2776 1559
rect 2832 1503 2859 1559
rect 2915 1503 2941 1559
rect 2997 1503 3009 1559
rect 2771 1498 3009 1503
use sky130_fd_io__gpio_ovtv2_hotswap_latch_i2c_fix  sky130_fd_io__gpio_ovtv2_hotswap_latch_i2c_fix_0
timestamp 1663361622
transform 1 0 -9399 0 1 -970
box 11695 1627 37770 16163
use sky130_fd_io__sio_hotswap_log_ovtv2_i2c_fix  sky130_fd_io__sio_hotswap_log_ovtv2_i2c_fix_0
timestamp 1663361622
transform 1 0 8920 0 1 1484
box 16 -95 6374 1336
<< labels >>
flabel metal1 s 12939 1513 12978 1541 0 FreeSans 200 0 0 0 EN_H
port 1 nsew
flabel metal1 s 12679 1475 12721 1503 0 FreeSans 200 0 0 0 FORCEHI_H[1]
port 2 nsew
flabel metal1 s 14236 1415 14338 1447 0 FreeSans 200 0 0 0 OD_I_H_N
port 3 nsew
flabel metal1 s 8613 1547 8663 1593 3 FreeSans 520 0 0 0 ENHS_LAT_H_N
port 4 nsew
flabel metal1 s 3224 2201 3334 2247 3 FreeSans 520 0 0 0 PGHS_H
port 5 nsew
flabel metal1 s 12400 1972 12429 2248 0 FreeSans 200 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 14371 1972 14400 2248 0 FreeSans 200 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 11555 1972 11581 2248 0 FreeSans 200 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 14371 2498 14400 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12400 2498 12429 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 14371 2424 14400 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12400 2424 12429 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 11522 2424 11542 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 11522 2498 11542 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12429 2424 12458 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12429 2498 12458 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 4800 823 5019 1016 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 5273 2579 5506 2710 3 FreeSans 520 0 0 0 VSSD
port 7 nsew
flabel metal1 s 3061 1511 3294 1626 3 FreeSans 520 0 0 0 VSSD
port 7 nsew
flabel metal1 s 9612 1287 9670 1329 0 FreeSans 440 0 0 0 VPWR_KA
port 8 nsew
flabel metal1 s 5354 1505 5412 1547 0 FreeSans 440 180 0 0 PAD_ESD
port 9 nsew
<< properties >>
string GDS_END 34147288
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 34132192
<< end >>
