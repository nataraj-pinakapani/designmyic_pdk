/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/xschem/decred_hash_macro/test2.spice