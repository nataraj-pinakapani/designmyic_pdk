magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 2 1 3 21 6 C0
port 1 nsew
rlabel  s 1 1 2 21 6 C0
port 1 nsew
rlabel  s 0 21 3 21 6 C0
port 1 nsew
rlabel  s 0 1 0 21 4 C0
port 1 nsew
rlabel  s 2 0 2 20 6 C1
port 2 nsew
rlabel  s 1 0 1 20 6 C1
port 2 nsew
rlabel  s 0 0 2 0 8 C1
port 2 nsew
rlabel metal_blue s 1 3 1 3 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 3 21
string LEFview TRUE
<< end >>
