magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel 
 s 1 13 25 16 6 VDDA
port 5 nsew power bidirectional
rlabel 
 s 51 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 13 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 51 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 75 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 75 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 14 75 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 14 75 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 13 75 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 13 75 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 14 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 14 74 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 13 74 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 13 74 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 16 74 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 15 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 14 74 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 14 74 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 13 74 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 74 13 74 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 14 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 14 73 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 13 73 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 13 73 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 14 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 14 73 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 13 73 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 73 13 73 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 73 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 14 73 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 14 73 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 13 73 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 13 73 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 14 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 14 72 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 13 72 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 13 72 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 16 72 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 15 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 14 72 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 14 72 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 13 72 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 72 13 72 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 14 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 14 71 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 13 71 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 13 71 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 14 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 14 71 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 13 71 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 71 13 71 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 71 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 14 71 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 14 71 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 13 71 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 13 71 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 14 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 14 70 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 13 70 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 13 70 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 16 70 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 15 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 14 70 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 14 70 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 13 70 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 70 13 70 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 14 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 14 69 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 13 69 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 13 69 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 16 69 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 15 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 14 69 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 14 69 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 13 69 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 69 13 69 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 14 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 14 68 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 13 68 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 13 68 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 14 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 14 68 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 13 68 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 68 13 68 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 68 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 14 68 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 14 68 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 13 68 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 13 68 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 14 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 14 67 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 13 67 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 13 67 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 16 67 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 15 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 14 67 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 14 67 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 13 67 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 67 13 67 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 14 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 14 66 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 13 66 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 13 66 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 14 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 14 66 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 13 66 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 66 13 66 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 66 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 14 66 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 14 66 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 13 66 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 13 66 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 14 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 14 65 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 13 65 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 13 65 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 16 65 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 15 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 14 65 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 14 65 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 13 65 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 65 13 65 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 14 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 14 64 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 13 64 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 13 64 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 14 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 14 64 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 13 64 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 64 13 64 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 64 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 14 64 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 14 64 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 13 64 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 13 64 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 14 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 14 63 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 13 63 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 13 63 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 16 63 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 15 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 14 63 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 14 63 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 13 63 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 63 13 63 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 14 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 14 62 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 13 62 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 13 62 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 14 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 14 62 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 13 62 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 62 13 62 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 62 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 14 62 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 14 62 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 13 62 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 13 62 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 14 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 14 61 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 13 61 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 13 61 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 16 61 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 15 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 14 61 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 14 61 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 13 61 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 61 13 61 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 14 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 14 60 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 13 60 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 13 60 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 14 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 14 60 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 13 60 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 60 13 60 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 60 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 14 60 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 14 60 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 13 60 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 13 60 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 14 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 14 59 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 13 59 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 13 59 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 16 59 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 15 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 14 59 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 14 59 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 13 59 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 59 13 59 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 14 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 14 58 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 13 58 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 13 58 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 14 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 14 58 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 13 58 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 58 13 58 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 58 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 14 58 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 14 58 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 13 58 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 13 58 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 14 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 14 57 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 13 57 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 13 57 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 16 57 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 15 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 14 57 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 14 57 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 13 57 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 57 13 57 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 14 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 14 56 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 13 56 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 13 56 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 14 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 14 56 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 13 56 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 56 13 56 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 56 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 14 56 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 14 56 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 13 56 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 13 56 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 14 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 14 55 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 13 55 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 13 55 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 16 55 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 15 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 14 55 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 14 55 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 13 55 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 55 13 55 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 14 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 14 54 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 13 54 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 13 54 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 14 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 14 54 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 13 54 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 54 13 54 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 54 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 14 54 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 14 54 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 13 54 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 13 54 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 16 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 15 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 14 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 14 53 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 13 53 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 53 13 53 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 53 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 14 53 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 14 53 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 13 53 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 13 53 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 14 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 14 52 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 13 52 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 13 52 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 16 52 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 15 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 14 52 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 14 52 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 13 52 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 52 13 52 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 14 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 14 51 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 13 51 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 13 51 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 16 51 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 15 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 14 51 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 14 51 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 13 51 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 51 13 51 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 14 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 14 24 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 13 24 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 13 24 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 14 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 14 24 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 13 24 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 24 13 24 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 24 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 14 24 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 14 24 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 13 24 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 13 24 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 14 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 14 23 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 13 23 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 13 23 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 16 23 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 15 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 14 23 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 14 23 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 13 23 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 23 13 23 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 14 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 14 22 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 13 22 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 13 22 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 14 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 14 22 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 13 22 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 22 13 22 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 22 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 14 22 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 14 22 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 13 22 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 13 22 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 14 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 14 21 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 13 21 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 13 21 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 16 21 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 15 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 14 21 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 14 21 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 13 21 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 21 13 21 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 14 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 14 20 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 13 20 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 13 20 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 14 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 14 20 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 13 20 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 20 13 20 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 20 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 14 20 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 14 20 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 13 20 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 13 20 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 14 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 14 19 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 13 19 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 13 19 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 16 19 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 15 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 14 19 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 14 19 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 13 19 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 19 13 19 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 14 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 14 18 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 13 18 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 13 18 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 14 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 14 18 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 13 18 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 18 13 18 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 18 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 14 18 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 14 18 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 13 18 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 13 18 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 14 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 14 17 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 13 17 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 13 17 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 16 17 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 15 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 14 17 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 14 17 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 13 17 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 17 13 17 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 14 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 14 16 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 13 16 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 13 16 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 14 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 14 16 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 13 16 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 16 13 16 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 16 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 14 16 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 14 16 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 13 16 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 13 16 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 16 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 15 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 14 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 14 15 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 13 15 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 15 13 15 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 15 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 14 15 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 14 15 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 13 15 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 13 15 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 14 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 14 14 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 13 14 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 13 14 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 16 14 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 15 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 14 14 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 14 14 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 13 14 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 14 13 14 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 14 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 14 13 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 13 13 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 13 13 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 14 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 14 13 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 13 13 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 13 13 13 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 13 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 14 13 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 14 13 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 13 13 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 13 13 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 14 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 14 12 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 13 12 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 13 12 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 16 12 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 15 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 14 12 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 14 12 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 13 12 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 12 13 12 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 14 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 14 11 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 13 11 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 13 11 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 14 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 14 11 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 13 11 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 11 13 11 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 11 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 14 11 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 14 11 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 13 11 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 13 11 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 14 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 14 10 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 13 10 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 13 10 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 16 10 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 15 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 14 10 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 14 10 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 13 10 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 10 13 10 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 14 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 14 9 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 13 9 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 13 9 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 14 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 14 9 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 13 9 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 9 13 9 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 9 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 14 9 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 14 9 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 13 9 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 13 9 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 14 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 14 8 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 13 8 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 13 8 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 16 8 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 15 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 14 8 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 14 8 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 13 8 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 8 13 8 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 14 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 14 7 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 13 7 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 13 7 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 14 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 14 7 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 13 7 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 7 13 7 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 7 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 14 7 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 14 7 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 13 7 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 13 7 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 14 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 14 6 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 13 6 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 13 6 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 16 6 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 15 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 14 6 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 14 6 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 13 6 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 6 13 6 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 14 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 14 5 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 13 5 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 13 5 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 14 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 14 5 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 13 5 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 5 13 5 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 5 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 14 5 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 14 5 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 13 5 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 13 5 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 14 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 14 4 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 13 4 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 13 4 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 16 4 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 15 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 14 4 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 14 4 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 13 4 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 4 13 4 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 14 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 14 3 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 13 3 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 13 3 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 14 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 14 3 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 13 3 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 3 13 3 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 3 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 14 3 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 14 3 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 13 3 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 13 3 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 14 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 14 2 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 13 2 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 13 2 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 16 2 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 15 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 14 2 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 14 2 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 13 2 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 2 13 2 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 14 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 14 1 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 13 1 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 13 1 13 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 16 1 16 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 15 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 14 1 15 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 14 1 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 13 1 14 6 VDDA
port 5 nsew power bidirectional
rlabel nfet_brown s 1 13 1 13 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 46 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 54 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 198
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
