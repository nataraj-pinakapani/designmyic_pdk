magic
tech minimum
timestamp 1644097874
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -7 -5 8 20
string LEFview TRUE
<< end >>
