magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1103 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 519 47 549 177
rect 603 47 633 177
rect 693 47 723 177
rect 777 47 807 177
rect 911 47 941 177
rect 995 47 1025 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 333 297 363 497
rect 421 297 451 497
rect 505 297 535 497
rect 693 297 723 497
rect 777 297 807 497
rect 911 297 941 497
rect 995 297 1025 497
<< ndiff >>
rect 27 101 79 177
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 101 247 177
rect 193 67 203 101
rect 237 67 247 101
rect 193 47 247 67
rect 277 95 331 177
rect 277 61 287 95
rect 321 61 331 95
rect 277 47 331 61
rect 361 165 413 177
rect 361 131 371 165
rect 405 131 413 165
rect 361 47 413 131
rect 467 165 519 177
rect 467 131 475 165
rect 509 131 519 165
rect 467 47 519 131
rect 549 95 603 177
rect 549 61 559 95
rect 593 61 603 95
rect 549 47 603 61
rect 633 101 693 177
rect 633 67 647 101
rect 681 67 693 101
rect 633 47 693 67
rect 723 93 777 177
rect 723 59 733 93
rect 767 59 777 93
rect 723 47 777 59
rect 807 101 911 177
rect 807 67 817 101
rect 851 67 911 101
rect 807 47 911 67
rect 941 93 995 177
rect 941 59 951 93
rect 985 59 995 93
rect 941 47 995 59
rect 1025 101 1077 177
rect 1025 67 1035 101
rect 1069 67 1077 101
rect 1025 47 1077 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 477 333 497
rect 277 443 287 477
rect 321 443 333 477
rect 277 409 333 443
rect 277 375 287 409
rect 321 375 333 409
rect 277 297 333 375
rect 363 485 421 497
rect 363 451 373 485
rect 407 451 421 485
rect 363 417 421 451
rect 363 383 373 417
rect 407 383 421 417
rect 363 297 421 383
rect 451 477 505 497
rect 451 443 461 477
rect 495 443 505 477
rect 451 409 505 443
rect 451 375 461 409
rect 495 375 505 409
rect 451 297 505 375
rect 535 485 587 497
rect 535 451 545 485
rect 579 451 587 485
rect 535 417 587 451
rect 535 383 545 417
rect 579 383 587 417
rect 535 297 587 383
rect 641 485 693 497
rect 641 451 649 485
rect 683 451 693 485
rect 641 297 693 451
rect 723 417 777 497
rect 723 383 733 417
rect 767 383 777 417
rect 723 349 777 383
rect 723 315 733 349
rect 767 315 777 349
rect 723 297 777 315
rect 807 485 911 497
rect 807 451 838 485
rect 872 451 911 485
rect 807 417 911 451
rect 807 383 838 417
rect 872 383 911 417
rect 807 297 911 383
rect 941 417 995 497
rect 941 383 951 417
rect 985 383 995 417
rect 941 349 995 383
rect 941 315 951 349
rect 985 315 995 349
rect 941 297 995 315
rect 1025 477 1077 497
rect 1025 443 1035 477
rect 1069 443 1077 477
rect 1025 409 1077 443
rect 1025 375 1035 409
rect 1069 375 1077 409
rect 1025 297 1077 375
<< ndiffc >>
rect 35 67 69 101
rect 119 59 153 93
rect 203 67 237 101
rect 287 61 321 95
rect 371 131 405 165
rect 475 131 509 165
rect 559 61 593 95
rect 647 67 681 101
rect 733 59 767 93
rect 817 67 851 101
rect 951 59 985 93
rect 1035 67 1069 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 443 153 477
rect 119 375 153 409
rect 203 451 237 485
rect 203 383 237 417
rect 287 443 321 477
rect 287 375 321 409
rect 373 451 407 485
rect 373 383 407 417
rect 461 443 495 477
rect 461 375 495 409
rect 545 451 579 485
rect 545 383 579 417
rect 649 451 683 485
rect 733 383 767 417
rect 733 315 767 349
rect 838 451 872 485
rect 838 383 872 417
rect 951 383 985 417
rect 951 315 985 349
rect 1035 443 1069 477
rect 1035 375 1069 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 333 497 363 523
rect 421 497 451 523
rect 505 497 535 523
rect 693 497 723 523
rect 777 497 807 523
rect 911 497 941 523
rect 995 497 1025 523
rect 79 265 109 297
rect 163 265 193 297
rect 22 249 193 265
rect 22 215 34 249
rect 68 215 102 249
rect 136 215 193 249
rect 22 199 193 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 265 277 297
rect 333 265 363 297
rect 421 265 451 297
rect 505 265 535 297
rect 693 265 723 297
rect 777 265 807 297
rect 247 249 369 265
rect 247 215 257 249
rect 291 215 325 249
rect 359 215 369 249
rect 247 199 369 215
rect 421 249 633 265
rect 421 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 633 249
rect 421 199 633 215
rect 683 249 807 265
rect 683 215 693 249
rect 727 215 761 249
rect 795 215 807 249
rect 683 199 807 215
rect 247 177 277 199
rect 331 177 361 199
rect 519 177 549 199
rect 603 177 633 199
rect 693 177 723 199
rect 777 177 807 199
rect 911 265 941 297
rect 995 265 1025 297
rect 911 261 1025 265
rect 911 249 1082 261
rect 911 215 964 249
rect 998 215 1032 249
rect 1066 215 1082 249
rect 911 203 1082 215
rect 911 199 1025 203
rect 911 177 941 199
rect 995 177 1025 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 519 21 549 47
rect 603 21 633 47
rect 693 21 723 47
rect 777 21 807 47
rect 911 21 941 47
rect 995 21 1025 47
<< polycont >>
rect 34 215 68 249
rect 102 215 136 249
rect 257 215 291 249
rect 325 215 359 249
rect 431 215 465 249
rect 499 215 533 249
rect 567 215 601 249
rect 693 215 727 249
rect 761 215 795 249
rect 964 215 998 249
rect 1032 215 1066 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 485 69 527
rect 19 451 35 485
rect 19 417 69 451
rect 19 383 35 417
rect 19 349 69 383
rect 19 315 35 349
rect 119 477 153 493
rect 119 409 153 443
rect 187 485 253 527
rect 187 451 203 485
rect 237 451 253 485
rect 187 417 253 451
rect 187 383 203 417
rect 237 383 253 417
rect 287 477 321 493
rect 287 409 321 443
rect 119 349 153 375
rect 357 485 427 527
rect 357 451 373 485
rect 407 451 427 485
rect 357 417 427 451
rect 357 383 373 417
rect 407 383 427 417
rect 461 477 495 493
rect 461 409 495 443
rect 287 349 321 375
rect 529 485 595 527
rect 822 485 888 493
rect 1035 485 1069 493
rect 529 451 545 485
rect 579 451 595 485
rect 629 451 649 485
rect 683 451 838 485
rect 872 477 1069 485
rect 872 451 1035 477
rect 529 417 595 451
rect 822 417 888 451
rect 529 383 545 417
rect 579 383 595 417
rect 717 383 733 417
rect 767 383 783 417
rect 822 383 838 417
rect 872 383 888 417
rect 932 383 951 417
rect 985 383 1001 417
rect 1035 409 1069 443
rect 461 349 495 375
rect 717 349 783 383
rect 119 315 733 349
rect 767 315 783 349
rect 932 349 998 383
rect 1035 359 1069 375
rect 932 336 951 349
rect 852 315 951 336
rect 985 315 1001 349
rect 19 299 69 315
rect 852 302 998 315
rect 27 249 160 265
rect 27 215 34 249
rect 68 215 102 249
rect 136 215 160 249
rect 27 199 160 215
rect 211 249 361 265
rect 211 215 257 249
rect 291 215 325 249
rect 359 215 361 249
rect 211 199 361 215
rect 400 249 623 265
rect 400 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 623 249
rect 400 199 623 215
rect 679 249 811 265
rect 679 215 693 249
rect 727 215 761 249
rect 795 215 811 249
rect 679 199 811 215
rect 852 165 895 302
rect 1035 259 1082 325
rect 946 249 1082 259
rect 946 215 964 249
rect 998 215 1032 249
rect 1066 215 1082 249
rect 35 131 371 165
rect 405 131 421 165
rect 459 131 475 165
rect 509 131 1069 165
rect 35 101 69 131
rect 203 101 237 131
rect 35 51 69 67
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 647 101 681 131
rect 203 51 237 67
rect 271 61 287 95
rect 321 61 559 95
rect 593 61 609 95
rect 817 101 851 131
rect 647 51 681 67
rect 717 59 733 93
rect 767 59 783 93
rect 717 17 783 59
rect 1035 101 1069 131
rect 817 51 851 67
rect 935 59 951 93
rect 985 59 1001 93
rect 935 17 1001 59
rect 1035 51 1069 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 948 221 982 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1040 221 1074 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 856 221 890 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 856 289 890 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 948 357 982 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 774 221 808 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1040 289 1074 323 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 494 221 528 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 856 153 890 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 682 221 716 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a311oi_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 3737180
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3726862
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 27.600 0.000 
<< end >>
