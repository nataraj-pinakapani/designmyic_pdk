magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 99 201 2483 203
rect 1 23 2483 201
rect 1 21 344 23
rect 610 21 1116 23
rect 2011 21 2483 23
rect 29 -17 63 21
<< scnmos >>
rect 80 47 110 175
rect 175 47 205 177
rect 404 49 434 177
rect 489 49 519 177
rect 691 47 721 175
rect 824 49 854 177
rect 1010 47 1040 177
rect 1112 49 1142 177
rect 1311 49 1341 177
rect 1396 49 1426 177
rect 1617 49 1647 177
rect 1705 49 1735 177
rect 1992 49 2022 177
rect 2087 47 2117 177
rect 2275 49 2305 177
rect 2370 47 2400 177
<< scpmoshvt >>
rect 80 297 110 497
rect 180 297 210 497
rect 404 297 434 465
rect 489 297 519 465
rect 702 297 732 465
rect 799 322 829 490
rect 1010 297 1040 497
rect 1112 297 1142 497
rect 1300 297 1330 465
rect 1384 297 1414 465
rect 1688 315 1718 483
rect 1772 315 1802 483
rect 1998 297 2028 497
rect 2082 297 2112 497
rect 2275 297 2305 497
rect 2359 297 2389 497
<< ndiff >>
rect 125 175 175 177
rect 27 161 80 175
rect 27 127 36 161
rect 70 127 80 161
rect 27 93 80 127
rect 27 59 36 93
rect 70 59 80 93
rect 27 47 80 59
rect 110 93 175 175
rect 110 59 126 93
rect 160 59 175 93
rect 110 47 175 59
rect 205 161 404 177
rect 205 127 215 161
rect 249 127 404 161
rect 205 93 404 127
rect 205 59 215 93
rect 249 59 360 93
rect 394 59 404 93
rect 205 49 404 59
rect 434 169 489 177
rect 434 135 444 169
rect 478 135 489 169
rect 434 49 489 135
rect 519 165 582 177
rect 758 175 824 177
rect 519 131 540 165
rect 574 131 582 165
rect 519 120 582 131
rect 519 49 581 120
rect 641 112 691 175
rect 636 101 691 112
rect 636 67 644 101
rect 678 67 691 101
rect 205 47 318 49
rect 636 47 691 67
rect 721 169 824 175
rect 721 135 780 169
rect 814 135 824 169
rect 721 49 824 135
rect 854 106 904 177
rect 958 165 1010 177
rect 958 131 966 165
rect 1000 131 1010 165
rect 958 121 1010 131
rect 959 120 1010 121
rect 854 105 905 106
rect 854 95 906 105
rect 854 61 864 95
rect 898 61 906 95
rect 854 49 906 61
rect 721 47 793 49
rect 960 47 1010 120
rect 1040 161 1112 177
rect 1040 127 1052 161
rect 1086 127 1112 161
rect 1040 93 1112 127
rect 1040 59 1052 93
rect 1086 59 1112 93
rect 1040 49 1112 59
rect 1142 133 1194 177
rect 1142 99 1152 133
rect 1186 99 1194 133
rect 1142 49 1194 99
rect 1251 114 1311 177
rect 1251 80 1267 114
rect 1301 80 1311 114
rect 1251 49 1311 80
rect 1341 169 1396 177
rect 1341 135 1351 169
rect 1385 135 1396 169
rect 1341 49 1396 135
rect 1426 169 1482 177
rect 1426 135 1436 169
rect 1470 135 1482 169
rect 1426 49 1482 135
rect 1565 122 1617 177
rect 1565 88 1573 122
rect 1607 88 1617 122
rect 1565 49 1617 88
rect 1647 169 1705 177
rect 1647 135 1661 169
rect 1695 135 1705 169
rect 1647 49 1705 135
rect 1735 153 1884 177
rect 1735 119 1761 153
rect 1795 119 1829 153
rect 1863 119 1884 153
rect 1735 49 1884 119
rect 1938 165 1992 177
rect 1938 131 1946 165
rect 1980 131 1992 165
rect 1938 97 1992 131
rect 1938 63 1946 97
rect 1980 63 1992 97
rect 1938 49 1992 63
rect 2022 97 2087 177
rect 2022 63 2036 97
rect 2070 63 2087 97
rect 2022 49 2087 63
rect 1040 47 1090 49
rect 2037 47 2087 49
rect 2117 165 2169 177
rect 2117 131 2127 165
rect 2161 131 2169 165
rect 2117 97 2169 131
rect 2117 63 2127 97
rect 2161 63 2169 97
rect 2117 47 2169 63
rect 2223 127 2275 177
rect 2223 93 2231 127
rect 2265 93 2275 127
rect 2223 49 2275 93
rect 2305 95 2370 177
rect 2305 61 2315 95
rect 2349 61 2370 95
rect 2305 49 2370 61
rect 2320 47 2370 49
rect 2400 163 2457 177
rect 2400 129 2415 163
rect 2449 129 2457 163
rect 2400 95 2457 129
rect 2400 61 2415 95
rect 2449 61 2457 95
rect 2400 47 2457 61
<< pdiff >>
rect 27 479 80 497
rect 27 445 36 479
rect 70 445 80 479
rect 27 411 80 445
rect 27 377 36 411
rect 70 377 80 411
rect 27 343 80 377
rect 27 309 36 343
rect 70 309 80 343
rect 27 297 80 309
rect 110 486 180 497
rect 110 452 120 486
rect 154 452 180 486
rect 110 297 180 452
rect 210 362 260 497
rect 633 493 683 505
rect 332 477 389 489
rect 332 443 344 477
rect 378 465 389 477
rect 378 443 404 465
rect 332 431 404 443
rect 210 350 298 362
rect 210 316 256 350
rect 290 316 298 350
rect 210 297 298 316
rect 354 297 404 431
rect 434 341 489 465
rect 434 307 444 341
rect 478 307 489 341
rect 434 297 489 307
rect 519 409 571 465
rect 519 375 529 409
rect 563 375 571 409
rect 519 297 571 375
rect 633 459 641 493
rect 675 465 683 493
rect 747 465 799 490
rect 675 459 702 465
rect 633 341 702 459
rect 633 307 658 341
rect 692 307 702 341
rect 633 297 702 307
rect 732 415 799 465
rect 732 381 742 415
rect 776 381 799 415
rect 732 322 799 381
rect 829 413 896 490
rect 829 379 839 413
rect 873 379 896 413
rect 829 322 896 379
rect 958 345 1010 497
rect 732 297 784 322
rect 958 311 966 345
rect 1000 311 1010 345
rect 958 297 1010 311
rect 1040 481 1112 497
rect 1040 447 1068 481
rect 1102 447 1112 481
rect 1040 297 1112 447
rect 1142 465 1269 497
rect 1904 483 1998 497
rect 1142 413 1300 465
rect 1142 379 1256 413
rect 1290 379 1300 413
rect 1142 345 1300 379
rect 1142 311 1152 345
rect 1186 311 1300 345
rect 1142 297 1300 311
rect 1330 341 1384 465
rect 1330 307 1340 341
rect 1374 307 1384 341
rect 1330 297 1384 307
rect 1414 409 1582 465
rect 1414 375 1476 409
rect 1510 375 1582 409
rect 1414 343 1582 375
rect 1636 441 1688 483
rect 1636 407 1644 441
rect 1678 407 1688 441
rect 1414 341 1580 343
rect 1414 307 1476 341
rect 1510 307 1580 341
rect 1636 315 1688 407
rect 1718 425 1772 483
rect 1718 391 1728 425
rect 1762 391 1772 425
rect 1718 357 1772 391
rect 1718 323 1728 357
rect 1762 323 1772 357
rect 1718 315 1772 323
rect 1802 341 1998 483
rect 1802 315 1952 341
rect 1414 297 1580 307
rect 1904 307 1952 315
rect 1986 307 1998 341
rect 1904 297 1998 307
rect 2028 489 2082 497
rect 2028 455 2038 489
rect 2072 455 2082 489
rect 2028 297 2082 455
rect 2112 479 2165 497
rect 2112 445 2123 479
rect 2157 445 2165 479
rect 2112 411 2165 445
rect 2112 377 2123 411
rect 2157 377 2165 411
rect 2112 343 2165 377
rect 2112 309 2123 343
rect 2157 309 2165 343
rect 2112 297 2165 309
rect 2223 480 2275 497
rect 2223 446 2231 480
rect 2265 446 2275 480
rect 2223 412 2275 446
rect 2223 378 2231 412
rect 2265 378 2275 412
rect 2223 344 2275 378
rect 2223 310 2231 344
rect 2265 310 2275 344
rect 2223 297 2275 310
rect 2305 475 2359 497
rect 2305 441 2315 475
rect 2349 441 2359 475
rect 2305 407 2359 441
rect 2305 373 2315 407
rect 2349 373 2359 407
rect 2305 297 2359 373
rect 2389 477 2446 497
rect 2389 443 2400 477
rect 2434 443 2446 477
rect 2389 409 2446 443
rect 2389 375 2400 409
rect 2434 375 2446 409
rect 2389 297 2446 375
<< ndiffc >>
rect 36 127 70 161
rect 36 59 70 93
rect 126 59 160 93
rect 215 127 249 161
rect 215 59 249 93
rect 360 59 394 93
rect 444 135 478 169
rect 540 131 574 165
rect 644 67 678 101
rect 780 135 814 169
rect 966 131 1000 165
rect 864 61 898 95
rect 1052 127 1086 161
rect 1052 59 1086 93
rect 1152 99 1186 133
rect 1267 80 1301 114
rect 1351 135 1385 169
rect 1436 135 1470 169
rect 1573 88 1607 122
rect 1661 135 1695 169
rect 1761 119 1795 153
rect 1829 119 1863 153
rect 1946 131 1980 165
rect 1946 63 1980 97
rect 2036 63 2070 97
rect 2127 131 2161 165
rect 2127 63 2161 97
rect 2231 93 2265 127
rect 2315 61 2349 95
rect 2415 129 2449 163
rect 2415 61 2449 95
<< pdiffc >>
rect 36 445 70 479
rect 36 377 70 411
rect 36 309 70 343
rect 120 452 154 486
rect 344 443 378 477
rect 256 316 290 350
rect 444 307 478 341
rect 529 375 563 409
rect 641 459 675 493
rect 658 307 692 341
rect 742 381 776 415
rect 839 379 873 413
rect 966 311 1000 345
rect 1068 447 1102 481
rect 1256 379 1290 413
rect 1152 311 1186 345
rect 1340 307 1374 341
rect 1476 375 1510 409
rect 1644 407 1678 441
rect 1476 307 1510 341
rect 1728 391 1762 425
rect 1728 323 1762 357
rect 1952 307 1986 341
rect 2038 455 2072 489
rect 2123 445 2157 479
rect 2123 377 2157 411
rect 2123 309 2157 343
rect 2231 446 2265 480
rect 2231 378 2265 412
rect 2231 310 2265 344
rect 2315 441 2349 475
rect 2315 373 2349 407
rect 2400 443 2434 477
rect 2400 375 2434 409
<< poly >>
rect 80 497 110 523
rect 180 497 210 523
rect 404 465 434 491
rect 489 465 519 491
rect 702 465 732 491
rect 799 490 829 516
rect 1010 497 1040 523
rect 1112 497 1142 523
rect 80 265 110 297
rect 180 265 210 297
rect 404 265 434 297
rect 67 249 133 265
rect 67 215 85 249
rect 119 215 133 249
rect 67 199 133 215
rect 175 249 262 265
rect 175 215 218 249
rect 252 215 262 249
rect 175 199 262 215
rect 304 249 434 265
rect 304 215 314 249
rect 348 215 434 249
rect 304 199 434 215
rect 80 175 110 199
rect 175 177 205 199
rect 404 177 434 199
rect 489 265 519 297
rect 702 265 732 297
rect 799 265 829 322
rect 1300 465 1330 491
rect 1384 465 1414 491
rect 1688 483 1718 509
rect 1772 483 1802 509
rect 1998 497 2028 523
rect 2082 497 2112 523
rect 2275 497 2305 523
rect 2359 497 2389 523
rect 1688 300 1718 315
rect 1010 265 1040 297
rect 1112 265 1142 297
rect 1300 265 1330 297
rect 1384 265 1414 297
rect 1599 270 1718 300
rect 1599 265 1647 270
rect 1772 265 1802 315
rect 1998 265 2028 297
rect 2082 265 2112 297
rect 2275 265 2305 297
rect 2359 265 2389 297
rect 489 249 732 265
rect 489 215 544 249
rect 578 215 732 249
rect 489 199 732 215
rect 797 249 1040 265
rect 797 215 848 249
rect 882 215 1040 249
rect 797 199 1040 215
rect 1082 249 1142 265
rect 1082 215 1092 249
rect 1126 215 1142 249
rect 1082 199 1142 215
rect 1241 249 1341 265
rect 1241 215 1251 249
rect 1285 215 1341 249
rect 1241 199 1341 215
rect 1384 249 1647 265
rect 1384 215 1573 249
rect 1607 215 1647 249
rect 1760 249 1814 265
rect 1760 222 1770 249
rect 1384 199 1647 215
rect 489 177 519 199
rect 691 175 721 199
rect 824 177 854 199
rect 1010 177 1040 199
rect 1112 177 1142 199
rect 1311 177 1341 199
rect 1396 177 1426 199
rect 1617 177 1647 199
rect 1705 215 1770 222
rect 1804 215 1814 249
rect 1705 199 1814 215
rect 1986 249 2040 265
rect 1986 215 1996 249
rect 2030 215 2040 249
rect 1986 199 2040 215
rect 2082 249 2305 265
rect 2082 215 2136 249
rect 2170 215 2305 249
rect 2082 199 2305 215
rect 2347 249 2401 265
rect 2347 215 2357 249
rect 2391 215 2401 249
rect 2347 199 2401 215
rect 1705 192 1811 199
rect 1705 177 1735 192
rect 1992 177 2022 199
rect 2087 177 2117 199
rect 2275 177 2305 199
rect 2370 177 2400 199
rect 80 21 110 47
rect 175 21 205 47
rect 404 21 434 49
rect 489 21 519 49
rect 691 21 721 47
rect 824 23 854 49
rect 1010 21 1040 47
rect 1112 23 1142 49
rect 1311 23 1341 49
rect 1396 23 1426 49
rect 1617 23 1647 49
rect 1705 21 1735 49
rect 1992 23 2022 49
rect 2087 21 2117 47
rect 2275 23 2305 49
rect 2370 21 2400 47
<< polycont >>
rect 85 215 119 249
rect 218 215 252 249
rect 314 215 348 249
rect 544 215 578 249
rect 848 215 882 249
rect 1092 215 1126 249
rect 1251 215 1285 249
rect 1573 215 1607 249
rect 1770 215 1804 249
rect 1996 215 2030 249
rect 2136 215 2170 249
rect 2357 215 2391 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 17 479 86 493
rect 17 445 36 479
rect 70 445 86 479
rect 17 411 86 445
rect 120 486 154 527
rect 343 477 641 493
rect 120 436 154 452
rect 188 443 344 477
rect 378 459 641 477
rect 675 459 703 493
rect 378 443 394 459
rect 17 377 36 411
rect 70 402 86 411
rect 188 402 222 443
rect 649 422 692 459
rect 70 377 222 402
rect 17 368 222 377
rect 256 391 290 409
rect 513 391 529 409
rect 17 343 88 368
rect 17 309 36 343
rect 70 309 88 343
rect 256 357 376 391
rect 513 357 514 391
rect 563 375 579 409
rect 548 357 579 375
rect 256 350 290 357
rect 17 300 88 309
rect 122 316 256 334
rect 122 300 290 316
rect 444 341 478 357
rect 658 341 692 422
rect 17 161 51 300
rect 122 265 156 300
rect 444 270 478 307
rect 85 249 156 265
rect 119 215 156 249
rect 190 249 268 255
rect 190 215 218 249
rect 252 215 268 249
rect 302 249 348 265
rect 302 215 314 249
rect 85 199 156 215
rect 122 181 156 199
rect 302 187 348 215
rect 122 161 265 181
rect 17 147 36 161
rect 20 127 36 147
rect 70 127 86 161
rect 122 147 215 161
rect 20 93 86 127
rect 199 127 215 147
rect 249 127 265 161
rect 302 153 305 187
rect 339 153 348 187
rect 302 133 348 153
rect 397 255 478 270
rect 431 221 478 255
rect 590 253 624 289
rect 560 249 624 253
rect 397 169 478 221
rect 528 215 544 249
rect 578 219 624 249
rect 578 215 594 219
rect 658 185 692 307
rect 742 458 1013 492
rect 742 415 776 458
rect 742 264 776 381
rect 816 413 889 424
rect 816 391 839 413
rect 816 357 828 391
rect 873 379 889 413
rect 963 413 1013 458
rect 1052 481 1118 527
rect 1052 447 1068 481
rect 1102 447 1118 481
rect 1165 459 1590 493
rect 1165 413 1199 459
rect 963 379 1199 413
rect 1240 413 1442 425
rect 1240 379 1256 413
rect 1290 391 1442 413
rect 1290 379 1306 391
rect 862 357 889 379
rect 816 339 889 357
rect 1240 345 1274 379
rect 938 323 966 345
rect 938 289 952 323
rect 1000 311 1034 345
rect 1127 311 1152 345
rect 1186 311 1274 345
rect 1340 341 1374 357
rect 986 289 1034 311
rect 938 277 1034 289
rect 966 265 1034 277
rect 742 230 814 264
rect 611 181 746 185
rect 397 135 444 169
rect 20 59 36 93
rect 70 59 86 93
rect 20 51 86 59
rect 126 93 160 109
rect 126 17 160 59
rect 199 93 265 127
rect 444 119 478 135
rect 524 165 746 181
rect 524 131 540 165
rect 574 151 746 165
rect 574 147 627 151
rect 574 131 605 147
rect 643 101 678 117
rect 643 93 644 101
rect 199 59 215 93
rect 249 59 360 93
rect 394 85 420 93
rect 503 85 644 93
rect 394 67 644 85
rect 394 59 678 67
rect 199 51 678 59
rect 712 85 746 151
rect 780 169 814 230
rect 780 119 814 135
rect 848 249 898 265
rect 882 215 898 249
rect 848 187 898 215
rect 848 153 857 187
rect 891 153 898 187
rect 848 129 898 153
rect 966 249 1126 265
rect 966 215 1092 249
rect 966 199 1126 215
rect 966 165 1000 199
rect 1160 163 1194 311
rect 1320 307 1340 335
rect 966 102 1000 131
rect 1036 127 1052 161
rect 1086 127 1102 161
rect 848 85 864 95
rect 712 61 864 85
rect 898 61 914 95
rect 712 51 914 61
rect 1036 93 1102 127
rect 1036 59 1052 93
rect 1086 59 1102 93
rect 1136 133 1194 163
rect 1228 255 1285 265
rect 1262 249 1285 255
rect 1228 215 1251 221
rect 1228 148 1285 215
rect 1320 185 1374 307
rect 1408 246 1442 391
rect 1476 409 1510 425
rect 1476 341 1510 375
rect 1556 344 1590 459
rect 1644 459 1882 493
rect 1644 441 1678 459
rect 1644 391 1678 407
rect 1712 391 1728 425
rect 1762 391 1778 425
rect 1712 357 1778 391
rect 1556 310 1607 344
rect 1476 306 1510 307
rect 1476 272 1522 306
rect 1488 258 1522 272
rect 1408 212 1454 246
rect 1488 221 1539 258
rect 1420 185 1454 212
rect 1504 187 1539 221
rect 1573 249 1607 310
rect 1573 199 1607 215
rect 1675 323 1728 357
rect 1762 323 1778 357
rect 1675 289 1688 323
rect 1722 306 1778 323
rect 1848 409 1882 459
rect 2038 489 2072 527
rect 2038 439 2072 455
rect 2107 479 2177 493
rect 2107 445 2123 479
rect 2157 445 2177 479
rect 2107 411 2177 445
rect 1848 408 2021 409
rect 1848 407 2024 408
rect 1848 406 2026 407
rect 1848 405 2029 406
rect 2107 405 2123 411
rect 1848 377 2123 405
rect 2157 377 2177 411
rect 1848 375 2177 377
rect 1722 289 1734 306
rect 1320 169 1385 185
rect 1320 151 1351 169
rect 1136 99 1152 133
rect 1186 99 1194 133
rect 1351 119 1385 135
rect 1420 169 1470 185
rect 1420 135 1436 169
rect 1420 119 1470 135
rect 1538 153 1539 187
rect 1675 185 1711 289
rect 1767 255 1814 265
rect 1767 249 1780 255
rect 1767 215 1770 249
rect 1804 215 1814 221
rect 1767 199 1814 215
rect 1136 76 1194 99
rect 1251 80 1267 114
rect 1301 85 1317 114
rect 1504 85 1539 153
rect 1661 169 1711 185
rect 1301 80 1539 85
rect 1036 17 1102 59
rect 1251 51 1539 80
rect 1573 122 1607 148
rect 1695 135 1711 169
rect 1848 153 1882 375
rect 2011 374 2177 375
rect 2014 373 2177 374
rect 2017 372 2177 373
rect 2020 371 2177 372
rect 2036 343 2177 371
rect 1661 119 1711 135
rect 1745 119 1761 153
rect 1795 119 1829 153
rect 1863 119 1882 153
rect 1928 307 1952 341
rect 1986 307 2002 341
rect 2036 309 2123 343
rect 2157 309 2177 343
rect 1928 165 1962 307
rect 2036 289 2177 309
rect 2215 480 2281 493
rect 2215 446 2231 480
rect 2265 446 2281 480
rect 2215 412 2281 446
rect 2215 378 2231 412
rect 2265 378 2281 412
rect 2215 344 2281 378
rect 2315 475 2366 527
rect 2349 441 2366 475
rect 2315 407 2366 441
rect 2349 373 2366 407
rect 2315 357 2366 373
rect 2400 477 2467 493
rect 2434 443 2467 477
rect 2400 409 2467 443
rect 2434 375 2467 409
rect 2400 357 2467 375
rect 2215 310 2231 344
rect 2265 310 2281 344
rect 2215 291 2281 310
rect 2036 265 2070 289
rect 1996 249 2070 265
rect 2030 215 2070 249
rect 2104 249 2193 255
rect 2104 215 2136 249
rect 2170 215 2193 249
rect 1996 199 2070 215
rect 2036 181 2070 199
rect 2231 187 2281 291
rect 2329 289 2336 323
rect 2370 289 2391 323
rect 2329 249 2391 289
rect 2329 215 2357 249
rect 2329 199 2391 215
rect 2036 165 2182 181
rect 1928 131 1946 165
rect 1980 131 1996 165
rect 2036 147 2127 165
rect 1573 85 1607 88
rect 1928 97 1996 131
rect 2106 131 2127 147
rect 2161 131 2182 165
rect 1928 85 1946 97
rect 1573 63 1946 85
rect 1980 63 1996 97
rect 1573 51 1996 63
rect 2036 97 2070 113
rect 2036 17 2070 63
rect 2106 97 2182 131
rect 2106 63 2127 97
rect 2161 63 2182 97
rect 2106 57 2182 63
rect 2231 153 2244 187
rect 2278 153 2281 187
rect 2425 165 2467 357
rect 2231 136 2281 153
rect 2399 163 2467 165
rect 2231 127 2265 136
rect 2399 129 2415 163
rect 2449 129 2467 163
rect 2231 54 2265 93
rect 2299 95 2365 102
rect 2299 61 2315 95
rect 2349 61 2365 95
rect 2299 17 2365 61
rect 2399 95 2467 129
rect 2399 61 2415 95
rect 2449 61 2467 95
rect 2399 51 2467 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 376 357 410 391
rect 514 375 529 391
rect 529 375 548 391
rect 514 357 548 375
rect 305 153 339 187
rect 397 221 431 255
rect 590 289 624 323
rect 828 379 839 391
rect 839 379 862 391
rect 828 357 862 379
rect 952 311 966 323
rect 966 311 986 323
rect 952 289 986 311
rect 857 153 891 187
rect 1228 249 1262 255
rect 1228 221 1251 249
rect 1251 221 1262 249
rect 1688 289 1722 323
rect 1504 153 1538 187
rect 1780 249 1814 255
rect 1780 221 1804 249
rect 1804 221 1814 249
rect 2336 289 2370 323
rect 2244 153 2278 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 364 391 422 397
rect 364 357 376 391
rect 410 388 422 391
rect 502 391 560 397
rect 502 388 514 391
rect 410 360 514 388
rect 410 357 422 360
rect 364 351 422 357
rect 502 357 514 360
rect 548 388 560 391
rect 816 391 874 397
rect 816 388 828 391
rect 548 360 828 388
rect 548 357 560 360
rect 502 351 560 357
rect 816 357 828 360
rect 862 357 874 391
rect 816 351 874 357
rect 578 323 636 329
rect 578 289 590 323
rect 624 320 636 323
rect 940 323 998 329
rect 940 320 952 323
rect 624 292 952 320
rect 624 289 636 292
rect 578 283 636 289
rect 940 289 952 292
rect 986 289 998 323
rect 940 283 998 289
rect 1676 323 1734 329
rect 1676 289 1688 323
rect 1722 320 1734 323
rect 2324 323 2382 329
rect 2324 320 2336 323
rect 1722 292 2336 320
rect 1722 289 1734 292
rect 1676 283 1734 289
rect 2324 289 2336 292
rect 2370 289 2382 323
rect 2324 283 2382 289
rect 385 255 443 261
rect 385 221 397 255
rect 431 252 443 255
rect 1216 255 1274 261
rect 1216 252 1228 255
rect 431 224 1228 252
rect 431 221 443 224
rect 385 215 443 221
rect 1216 221 1228 224
rect 1262 252 1274 255
rect 1768 255 1826 261
rect 1768 252 1780 255
rect 1262 224 1780 252
rect 1262 221 1274 224
rect 1216 215 1274 221
rect 1768 221 1780 224
rect 1814 221 1826 255
rect 1768 215 1826 221
rect 293 187 351 193
rect 293 153 305 187
rect 339 184 351 187
rect 845 187 903 193
rect 845 184 857 187
rect 339 156 857 184
rect 339 153 351 156
rect 293 147 351 153
rect 845 153 857 156
rect 891 153 903 187
rect 845 147 903 153
rect 1492 187 1550 193
rect 1492 153 1504 187
rect 1538 184 1550 187
rect 2232 187 2290 193
rect 2232 184 2244 187
rect 1538 156 2244 184
rect 1538 153 1550 156
rect 1492 147 1550 153
rect 2232 153 2244 156
rect 2278 153 2290 187
rect 2232 147 2290 153
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
flabel locali s 1320 289 1354 323 0 FreeSans 300 0 0 0 COUT
port 8 nsew signal output
flabel locali s 305 153 339 187 0 FreeSans 300 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 300 180 0 0 A
port 1 nsew signal input
flabel locali s 2428 221 2462 255 0 FreeSans 300 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2148 221 2182 255 0 FreeSans 300 0 0 0 CIN
port 3 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 322 170 322 170 0 FreeSans 300 0 0 0 B
port 2 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fahcin_1
rlabel locali s 848 129 898 265 1 B
port 2 nsew signal input
rlabel metal1 s 845 184 903 193 1 B
port 2 nsew signal input
rlabel metal1 s 845 147 903 156 1 B
port 2 nsew signal input
rlabel metal1 s 293 184 351 193 1 B
port 2 nsew signal input
rlabel metal1 s 293 156 903 184 1 B
port 2 nsew signal input
rlabel metal1 s 293 147 351 156 1 B
port 2 nsew signal input
rlabel metal1 s 0 -48 2484 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2484 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2484 544
string GDS_END 2132810
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 2113526
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 62.100 13.600 
<< end >>
