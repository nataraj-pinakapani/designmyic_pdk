/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/sky130_fd_pr__diode_pd2nw_05v5_lvt_fail.cdl