magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 4 43 998 283
rect -26 -43 1082 43
<< locali >>
rect 112 355 302 411
rect 409 355 647 430
rect 268 319 302 355
rect 683 319 743 367
rect 268 301 743 319
rect 268 285 717 301
rect 793 265 874 485
rect 770 99 874 265
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 26 521 76 751
rect 112 735 506 751
rect 146 701 184 735
rect 218 701 256 735
rect 290 701 328 735
rect 362 701 400 735
rect 434 701 472 735
rect 112 557 506 701
rect 542 625 576 751
rect 612 735 944 751
rect 612 701 617 735
rect 651 701 689 735
rect 723 701 761 735
rect 795 701 833 735
rect 867 701 905 735
rect 939 701 944 735
rect 612 661 944 701
rect 980 625 1030 751
rect 542 591 1030 625
rect 542 557 576 591
rect 612 521 944 555
rect 26 487 646 521
rect 26 319 76 487
rect 26 285 232 319
rect 18 113 136 249
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 136 113
rect 182 99 232 285
rect 910 399 944 521
rect 980 435 1030 591
rect 910 333 976 399
rect 268 113 734 249
rect 18 73 136 79
rect 302 79 340 113
rect 374 79 412 113
rect 446 79 484 113
rect 518 79 556 113
rect 590 79 628 113
rect 662 79 700 113
rect 910 113 1028 265
rect 268 73 734 79
rect 910 79 916 113
rect 950 79 988 113
rect 1022 79 1028 113
rect 910 73 1028 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 112 701 146 735
rect 184 701 218 735
rect 256 701 290 735
rect 328 701 362 735
rect 400 701 434 735
rect 472 701 506 735
rect 617 701 651 735
rect 689 701 723 735
rect 761 701 795 735
rect 833 701 867 735
rect 905 701 939 735
rect 24 79 58 113
rect 96 79 130 113
rect 268 79 302 113
rect 340 79 374 113
rect 412 79 446 113
rect 484 79 518 113
rect 556 79 590 113
rect 628 79 662 113
rect 700 79 734 113
rect 916 79 950 113
rect 988 79 1022 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 735 1056 763
rect 0 701 112 735
rect 146 701 184 735
rect 218 701 256 735
rect 290 701 328 735
rect 362 701 400 735
rect 434 701 472 735
rect 506 701 617 735
rect 651 701 689 735
rect 723 701 761 735
rect 795 701 833 735
rect 867 701 905 735
rect 939 701 1056 735
rect 0 689 1056 701
rect 0 113 1056 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 268 113
rect 302 79 340 113
rect 374 79 412 113
rect 446 79 484 113
rect 518 79 556 113
rect 590 79 628 113
rect 662 79 700 113
rect 734 79 916 113
rect 950 79 988 113
rect 1022 79 1056 113
rect 0 51 1056 79
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel locali s 409 355 647 430 6 A
port 1 nsew signal input
rlabel locali s 268 285 717 301 6 B
port 2 nsew signal input
rlabel locali s 268 301 743 319 6 B
port 2 nsew signal input
rlabel locali s 683 319 743 367 6 B
port 2 nsew signal input
rlabel locali s 268 319 302 355 6 B
port 2 nsew signal input
rlabel locali s 112 355 302 411 6 B
port 2 nsew signal input
rlabel metal1 s 0 51 1056 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 1056 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 1082 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 43 998 283 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 1056 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 1122 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 1056 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 770 99 874 265 6 X
port 7 nsew signal output
rlabel locali s 793 265 874 485 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1056 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 743414
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 731354
<< end >>
