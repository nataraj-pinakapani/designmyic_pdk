magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 64 36 67 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel  s 39 64 80 67 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel  s 0 59 52 62 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel  s 54 59 80 62 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel � s 51 0 51 2 6 ANALOG_EN
port 22 nsew signal input
rlabel � s 44 0 45 2 6 ANALOG_POL
port 26 nsew signal input
rlabel � s 29 0 29 2 6 ANALOG_SEL
port 23 nsew signal input
rlabel � s 26 0 26 2 6 DM[2]
port 6 nsew signal input
rlabel � s 57 0 57 2 6 DM[1]
port 7 nsew signal input
rlabel � s 47 0 48 2 6 DM[0]
port 8 nsew signal input
rlabel � s 35 0 35 2 6 ENABLE_H
port 13 nsew signal input
rlabel � s 38 0 39 2 6 ENABLE_INP_H
port 15 nsew signal input
rlabel � s 13 0 14 2 6 ENABLE_VDDA_H
port 14 nsew signal input
rlabel � s 69 0 69 2 6 ENABLE_VDDIO
port 24 nsew signal input
rlabel � s 17 0 17 2 6 ENABLE_VSWITCH_H
port 25 nsew signal input
rlabel � s 32 0 32 2 6 HLD_H_N
port 9 nsew signal input
rlabel � s 23 0 23 2 6 HLD_OVR
port 21 nsew signal input
rlabel � s 7 0 8 2 6 IB_MODE_SEL
port 12 nsew signal input
rlabel � s 75 0 75 2 6 IN
port 10 nsew signal output
rlabel � s 1 0 2 2 6 IN_H
port 1 nsew signal output
rlabel � s 42 0 42 2 6 INP_DIS
port 11 nsew signal input
rlabel � s 4 0 5 2 6 OE_N
port 16 nsew signal input
rlabel � s 20 0 20 2 6 OUT
port 27 nsew signal input
rlabel  s 11 116 74 178 6 PAD
port 5 nsew signal bidirectional
rlabel � s 63 0 63 2 6 PAD_A_ESD_0_H
port 3 nsew signal bidirectional
rlabel � s 60 0 60 2 6 PAD_A_ESD_1_H
port 4 nsew signal bidirectional
rlabel � s 53 0 54 2 6 PAD_A_NOESD_H
port 2 nsew signal bidirectional
rlabel � s 66 0 66 2 6 SLOW
port 19 nsew signal input
rlabel � s 72 0 72 2 6 TIE_HI_ESD
port 17 nsew signal output
rlabel � s 78 0 79 2 6 TIE_LO_ESD
port 18 nsew signal output
rlabel  s 0 20 1 24 4 VCCD
port 36 nsew power bidirectional
rlabel  s 0 20 1 25 4 VCCD
port 36 nsew power bidirectional
rlabel  s 79 20 80 24 6 VCCD
port 36 nsew power bidirectional
rlabel  s 79 20 80 25 6 VCCD
port 36 nsew power bidirectional
rlabel  s 0 13 1 18 4 VCCHIB
port 34 nsew power bidirectional
rlabel  s 0 13 1 18 4 VCCHIB
port 34 nsew power bidirectional
rlabel  s 79 13 80 18 6 VCCHIB
port 34 nsew power bidirectional
rlabel  s 79 13 80 18 6 VCCHIB
port 34 nsew power bidirectional
rlabel  s 0 26 1 29 4 VDDA
port 31 nsew power bidirectional
rlabel  s 0 26 1 29 4 VDDA
port 31 nsew power bidirectional
rlabel  s 79 26 80 29 6 VDDA
port 31 nsew power bidirectional
rlabel  s 79 26 80 29 6 VDDA
port 31 nsew power bidirectional
rlabel  s 0 81 1 106 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 31 1 35 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 31 1 35 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 81 1 106 4 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 81 80 106 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 31 80 35 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 31 80 35 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 79 81 80 106 6 VDDIO
port 35 nsew power bidirectional
rlabel  s 0 75 1 79 4 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 0 75 1 80 4 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 79 75 80 79 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 79 75 80 80 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel  s 0 59 1 68 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 48 1 51 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 59 3 59 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 63 1 64 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 67 3 68 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 48 1 51 4 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 59 80 68 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 48 80 51 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 63 80 64 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 47 67 80 68 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 47 59 80 59 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 79 48 80 51 6 VSSA
port 30 nsew ground bidirectional
rlabel  s 0 53 1 57 4 VSSD
port 38 nsew ground bidirectional
rlabel  s 0 53 1 57 4 VSSD
port 38 nsew ground bidirectional
rlabel  s 79 53 80 57 6 VSSD
port 38 nsew ground bidirectional
rlabel  s 79 53 80 57 6 VSSD
port 38 nsew ground bidirectional
rlabel  s 0 187 1 211 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 37 1 41 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 37 1 41 4 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 187 80 211 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 37 80 41 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 79 37 80 41 6 VSSIO
port 37 nsew ground bidirectional
rlabel  s 0 69 1 74 4 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 0 69 1 74 4 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 79 69 80 74 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 79 69 80 74 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel  s 0 43 1 46 4 VSWITCH
port 32 nsew power bidirectional
rlabel  s 0 43 1 46 4 VSWITCH
port 32 nsew power bidirectional
rlabel  s 79 43 80 46 6 VSWITCH
port 32 nsew power bidirectional
rlabel  s 79 43 80 46 6 VSWITCH
port 32 nsew power bidirectional
rlabel � s 11 0 11 2 6 VTRIP_SEL
port 20 nsew signal input
<< properties >>
string LEFclass PAD INOUT
string FIXED_BBOX 0 0 80 211
string LEFview TRUE
<< end >>
