magic
tech minimum
timestamp 1644097874
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -91 -91 93 91
string LEFview TRUE
string gencell sky130_fd_pr__rf_test_coil3
string library sky130
string parameter m=1
<< end >>
