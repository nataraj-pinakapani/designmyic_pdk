magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 5190 2009 5884 2225
rect 13942 1725 14274 2219
<< pwell >>
rect 89 2703 741 2716
rect 89 2289 1123 2703
rect 89 1740 741 2289
rect 89 1407 849 1740
rect 89 1398 741 1407
<< mvnmos >>
rect 115 2537 715 2637
rect 897 2524 1097 2624
rect 897 2368 1097 2468
rect 115 2257 715 2357
rect 115 2101 715 2201
rect 115 1945 715 2045
rect 115 1789 715 1889
rect 115 1633 715 1733
rect 115 1477 715 1577
<< mvpmos >>
rect 5309 2075 5509 2159
rect 5565 2075 5765 2159
rect 14008 2000 14208 2100
rect 14008 1844 14208 1944
<< mvndiff >>
rect 115 2682 715 2690
rect 115 2648 193 2682
rect 227 2648 261 2682
rect 295 2648 329 2682
rect 363 2648 397 2682
rect 431 2648 465 2682
rect 499 2648 533 2682
rect 567 2648 601 2682
rect 635 2648 669 2682
rect 703 2648 715 2682
rect 115 2637 715 2648
rect 897 2669 1097 2677
rect 897 2635 909 2669
rect 943 2635 977 2669
rect 1011 2635 1045 2669
rect 1079 2635 1097 2669
rect 897 2624 1097 2635
rect 115 2526 715 2537
rect 115 2492 193 2526
rect 227 2492 261 2526
rect 295 2492 329 2526
rect 363 2492 397 2526
rect 431 2492 465 2526
rect 499 2492 533 2526
rect 567 2492 601 2526
rect 635 2492 669 2526
rect 703 2492 715 2526
rect 115 2484 715 2492
rect 897 2513 1097 2524
rect 897 2479 909 2513
rect 943 2479 977 2513
rect 1011 2479 1045 2513
rect 1079 2479 1097 2513
rect 897 2468 1097 2479
rect 115 2402 715 2410
rect 115 2368 193 2402
rect 227 2368 261 2402
rect 295 2368 329 2402
rect 363 2368 397 2402
rect 431 2368 465 2402
rect 499 2368 533 2402
rect 567 2368 601 2402
rect 635 2368 669 2402
rect 703 2368 715 2402
rect 115 2357 715 2368
rect 897 2357 1097 2368
rect 897 2323 909 2357
rect 943 2323 977 2357
rect 1011 2323 1045 2357
rect 1079 2323 1097 2357
rect 897 2315 1097 2323
rect 115 2246 715 2257
rect 115 2212 193 2246
rect 227 2212 261 2246
rect 295 2212 329 2246
rect 363 2212 397 2246
rect 431 2212 465 2246
rect 499 2212 533 2246
rect 567 2212 601 2246
rect 635 2212 669 2246
rect 703 2212 715 2246
rect 115 2201 715 2212
rect 115 2090 715 2101
rect 115 2056 193 2090
rect 227 2056 261 2090
rect 295 2056 329 2090
rect 363 2056 397 2090
rect 431 2056 465 2090
rect 499 2056 533 2090
rect 567 2056 601 2090
rect 635 2056 669 2090
rect 703 2056 715 2090
rect 115 2045 715 2056
rect 115 1934 715 1945
rect 115 1900 193 1934
rect 227 1900 261 1934
rect 295 1900 329 1934
rect 363 1900 397 1934
rect 431 1900 465 1934
rect 499 1900 533 1934
rect 567 1900 601 1934
rect 635 1900 669 1934
rect 703 1900 715 1934
rect 115 1889 715 1900
rect 115 1778 715 1789
rect 115 1744 193 1778
rect 227 1744 261 1778
rect 295 1744 329 1778
rect 363 1744 397 1778
rect 431 1744 465 1778
rect 499 1744 533 1778
rect 567 1744 601 1778
rect 635 1744 669 1778
rect 703 1744 715 1778
rect 115 1733 715 1744
rect 115 1622 715 1633
rect 115 1588 193 1622
rect 227 1588 261 1622
rect 295 1588 329 1622
rect 363 1588 397 1622
rect 431 1588 465 1622
rect 499 1588 533 1622
rect 567 1588 601 1622
rect 635 1588 669 1622
rect 703 1588 715 1622
rect 115 1577 715 1588
rect 115 1466 715 1477
rect 115 1432 193 1466
rect 227 1432 261 1466
rect 295 1432 329 1466
rect 363 1432 397 1466
rect 431 1432 465 1466
rect 499 1432 533 1466
rect 567 1432 601 1466
rect 635 1432 669 1466
rect 703 1432 715 1466
rect 115 1424 715 1432
<< mvpdiff >>
rect 5256 2147 5309 2159
rect 5256 2113 5264 2147
rect 5298 2113 5309 2147
rect 5256 2075 5309 2113
rect 5509 2147 5565 2159
rect 5509 2113 5520 2147
rect 5554 2113 5565 2147
rect 5509 2075 5565 2113
rect 5765 2147 5818 2159
rect 5765 2113 5776 2147
rect 5810 2113 5818 2147
rect 5765 2075 5818 2113
rect 14008 2145 14208 2153
rect 14008 2111 14020 2145
rect 14054 2111 14088 2145
rect 14122 2111 14156 2145
rect 14190 2111 14208 2145
rect 14008 2100 14208 2111
rect 14008 1989 14208 2000
rect 14008 1955 14020 1989
rect 14054 1955 14088 1989
rect 14122 1955 14156 1989
rect 14190 1955 14208 1989
rect 14008 1944 14208 1955
rect 14008 1833 14208 1844
rect 14008 1799 14020 1833
rect 14054 1799 14088 1833
rect 14122 1799 14156 1833
rect 14190 1799 14208 1833
rect 14008 1791 14208 1799
<< mvndiffc >>
rect 193 2648 227 2682
rect 261 2648 295 2682
rect 329 2648 363 2682
rect 397 2648 431 2682
rect 465 2648 499 2682
rect 533 2648 567 2682
rect 601 2648 635 2682
rect 669 2648 703 2682
rect 909 2635 943 2669
rect 977 2635 1011 2669
rect 1045 2635 1079 2669
rect 193 2492 227 2526
rect 261 2492 295 2526
rect 329 2492 363 2526
rect 397 2492 431 2526
rect 465 2492 499 2526
rect 533 2492 567 2526
rect 601 2492 635 2526
rect 669 2492 703 2526
rect 909 2479 943 2513
rect 977 2479 1011 2513
rect 1045 2479 1079 2513
rect 193 2368 227 2402
rect 261 2368 295 2402
rect 329 2368 363 2402
rect 397 2368 431 2402
rect 465 2368 499 2402
rect 533 2368 567 2402
rect 601 2368 635 2402
rect 669 2368 703 2402
rect 909 2323 943 2357
rect 977 2323 1011 2357
rect 1045 2323 1079 2357
rect 193 2212 227 2246
rect 261 2212 295 2246
rect 329 2212 363 2246
rect 397 2212 431 2246
rect 465 2212 499 2246
rect 533 2212 567 2246
rect 601 2212 635 2246
rect 669 2212 703 2246
rect 193 2056 227 2090
rect 261 2056 295 2090
rect 329 2056 363 2090
rect 397 2056 431 2090
rect 465 2056 499 2090
rect 533 2056 567 2090
rect 601 2056 635 2090
rect 669 2056 703 2090
rect 193 1900 227 1934
rect 261 1900 295 1934
rect 329 1900 363 1934
rect 397 1900 431 1934
rect 465 1900 499 1934
rect 533 1900 567 1934
rect 601 1900 635 1934
rect 669 1900 703 1934
rect 193 1744 227 1778
rect 261 1744 295 1778
rect 329 1744 363 1778
rect 397 1744 431 1778
rect 465 1744 499 1778
rect 533 1744 567 1778
rect 601 1744 635 1778
rect 669 1744 703 1778
rect 193 1588 227 1622
rect 261 1588 295 1622
rect 329 1588 363 1622
rect 397 1588 431 1622
rect 465 1588 499 1622
rect 533 1588 567 1622
rect 601 1588 635 1622
rect 669 1588 703 1622
rect 193 1432 227 1466
rect 261 1432 295 1466
rect 329 1432 363 1466
rect 397 1432 431 1466
rect 465 1432 499 1466
rect 533 1432 567 1466
rect 601 1432 635 1466
rect 669 1432 703 1466
<< mvpdiffc >>
rect 5264 2113 5298 2147
rect 5520 2113 5554 2147
rect 5776 2113 5810 2147
rect 14020 2111 14054 2145
rect 14088 2111 14122 2145
rect 14156 2111 14190 2145
rect 14020 1955 14054 1989
rect 14088 1955 14122 1989
rect 14156 1955 14190 1989
rect 14020 1799 14054 1833
rect 14088 1799 14122 1833
rect 14156 1799 14190 1833
<< psubdiff >>
rect 789 1690 823 1714
rect 789 1591 823 1656
rect 789 1491 823 1557
rect 789 1433 823 1457
<< psubdiffcont >>
rect 789 1656 823 1690
rect 789 1557 823 1591
rect 789 1457 823 1491
<< poly >>
rect 17 2638 83 2654
rect 17 2604 33 2638
rect 67 2637 83 2638
rect 67 2604 115 2637
rect 17 2570 115 2604
rect 17 2536 33 2570
rect 67 2537 115 2570
rect 715 2537 747 2637
rect 1127 2645 1193 2661
rect 1127 2624 1143 2645
rect 67 2536 83 2537
rect 17 2520 83 2536
rect 865 2524 897 2624
rect 1097 2611 1143 2624
rect 1177 2611 1193 2645
rect 1097 2574 1193 2611
rect 1097 2540 1143 2574
rect 1177 2540 1193 2574
rect 1097 2524 1193 2540
rect 865 2368 897 2468
rect 1097 2452 1193 2468
rect 1097 2418 1143 2452
rect 1177 2418 1193 2452
rect 1097 2381 1193 2418
rect 1097 2368 1143 2381
rect 17 2341 115 2357
rect 17 2307 33 2341
rect 67 2307 115 2341
rect 17 2271 115 2307
rect 17 2237 33 2271
rect 67 2257 115 2271
rect 715 2257 747 2357
rect 1127 2347 1143 2368
rect 1177 2347 1193 2381
rect 1127 2331 1193 2347
rect 67 2237 83 2257
rect 17 2202 83 2237
rect 17 2168 33 2202
rect 67 2201 83 2202
rect 5309 2241 5509 2257
rect 5309 2207 5325 2241
rect 5359 2207 5459 2241
rect 5493 2207 5509 2241
rect 67 2168 115 2201
rect 17 2133 115 2168
rect 17 2099 33 2133
rect 67 2101 115 2133
rect 715 2101 747 2201
rect 5309 2159 5509 2207
rect 5565 2241 5765 2257
rect 5565 2207 5581 2241
rect 5615 2207 5715 2241
rect 5749 2207 5765 2241
rect 5565 2159 5765 2207
rect 67 2099 83 2101
rect 17 2064 83 2099
rect 17 2030 33 2064
rect 67 2045 83 2064
rect 67 2030 115 2045
rect 17 1995 115 2030
rect 17 1961 33 1995
rect 67 1961 115 1995
rect 17 1945 115 1961
rect 715 1945 747 2045
rect 5309 2043 5509 2075
rect 5565 2043 5765 2075
rect 13976 2000 14008 2100
rect 14208 2084 14306 2100
rect 14208 2050 14256 2084
rect 14290 2050 14306 2084
rect 14208 2000 14306 2050
rect 14240 1989 14306 2000
rect 14240 1955 14256 1989
rect 14290 1955 14306 1989
rect 14240 1944 14306 1955
rect 17 1873 115 1889
rect 17 1839 33 1873
rect 67 1839 115 1873
rect 17 1803 115 1839
rect 17 1769 33 1803
rect 67 1789 115 1803
rect 715 1789 747 1889
rect 13976 1844 14008 1944
rect 14208 1894 14306 1944
rect 14208 1860 14256 1894
rect 14290 1860 14306 1894
rect 14208 1844 14306 1860
rect 67 1769 83 1789
rect 17 1734 83 1769
rect 17 1700 33 1734
rect 67 1733 83 1734
rect 67 1700 115 1733
rect 17 1665 115 1700
rect 17 1631 33 1665
rect 67 1633 115 1665
rect 715 1633 747 1733
rect 67 1631 83 1633
rect 17 1596 83 1631
rect 17 1562 33 1596
rect 67 1577 83 1596
rect 67 1562 115 1577
rect 17 1527 115 1562
rect 17 1493 33 1527
rect 67 1493 115 1527
rect 17 1477 115 1493
rect 715 1477 747 1577
<< polycont >>
rect 33 2604 67 2638
rect 33 2536 67 2570
rect 1143 2611 1177 2645
rect 1143 2540 1177 2574
rect 1143 2418 1177 2452
rect 33 2307 67 2341
rect 33 2237 67 2271
rect 1143 2347 1177 2381
rect 33 2168 67 2202
rect 5325 2207 5359 2241
rect 5459 2207 5493 2241
rect 33 2099 67 2133
rect 5581 2207 5615 2241
rect 5715 2207 5749 2241
rect 33 2030 67 2064
rect 33 1961 67 1995
rect 14256 2050 14290 2084
rect 14256 1955 14290 1989
rect 33 1839 67 1873
rect 33 1769 67 1803
rect 14256 1860 14290 1894
rect 33 1700 67 1734
rect 33 1631 67 1665
rect 33 1562 67 1596
rect 33 1493 67 1527
<< locali >>
rect -31 2642 67 2654
rect 177 2648 193 2682
rect 227 2648 261 2682
rect 295 2648 329 2682
rect 363 2648 397 2682
rect 431 2648 465 2682
rect 499 2648 531 2682
rect 567 2648 601 2682
rect 635 2648 669 2682
rect 707 2648 719 2682
rect -3 2638 67 2642
rect -3 2608 33 2638
rect -37 2604 33 2608
rect -37 2570 67 2604
rect -37 2566 33 2570
rect -3 2536 33 2566
rect -3 2532 67 2536
rect -31 2520 67 2532
rect 793 2613 827 2654
rect 893 2635 909 2669
rect 943 2635 977 2669
rect 1011 2635 1045 2669
rect 1083 2635 1095 2669
rect 1143 2649 1177 2661
rect 793 2538 827 2579
rect 177 2492 193 2526
rect 227 2492 261 2526
rect 295 2492 329 2526
rect 363 2492 397 2526
rect 431 2492 465 2526
rect 499 2492 531 2526
rect 567 2492 601 2526
rect 637 2492 669 2526
rect 703 2492 719 2526
rect 1143 2574 1177 2611
rect 1143 2524 1177 2536
rect 793 2463 827 2504
rect 903 2479 909 2513
rect 975 2479 977 2513
rect 1011 2479 1045 2513
rect 1079 2479 1095 2513
rect 177 2368 193 2402
rect 227 2368 261 2402
rect 322 2368 329 2402
rect 394 2368 397 2402
rect 431 2368 465 2402
rect 499 2368 533 2402
rect 567 2368 601 2402
rect 635 2368 669 2402
rect 703 2368 719 2402
rect 793 2388 827 2429
rect 33 2345 67 2357
rect 64 2341 67 2345
rect 30 2307 33 2311
rect 30 2271 67 2307
rect 30 2256 33 2271
rect 1143 2456 1177 2468
rect 1143 2381 1177 2418
rect 793 2313 827 2354
rect 893 2323 909 2357
rect 943 2323 977 2357
rect 1011 2323 1045 2357
rect 1083 2323 1095 2357
rect 1143 2331 1177 2343
rect 64 2222 67 2237
rect 30 2202 67 2222
rect 177 2212 193 2246
rect 227 2212 261 2246
rect 295 2212 329 2246
rect 363 2212 397 2246
rect 431 2212 465 2246
rect 499 2212 531 2246
rect 567 2212 601 2246
rect 637 2212 669 2246
rect 703 2212 719 2246
rect 793 2238 827 2279
rect 30 2168 33 2202
rect 30 2167 67 2168
rect 64 2133 67 2167
rect 30 2099 33 2133
rect 30 2079 67 2099
rect 793 2163 827 2204
rect 64 2064 67 2079
rect 177 2056 193 2090
rect 227 2056 261 2090
rect 322 2056 329 2090
rect 394 2056 397 2090
rect 431 2056 465 2090
rect 499 2056 533 2090
rect 567 2056 601 2090
rect 635 2056 669 2090
rect 703 2056 719 2090
rect 793 2087 827 2129
rect 5154 2211 5231 2245
rect 5612 2241 5680 2248
rect 5154 2163 5265 2211
rect 5309 2207 5325 2241
rect 5359 2207 5459 2241
rect 5493 2207 5509 2241
rect 5565 2214 5578 2241
rect 5615 2214 5680 2241
rect 5714 2214 5715 2241
rect 5565 2207 5581 2214
rect 5615 2207 5715 2214
rect 5749 2207 5765 2241
rect 5364 2167 5470 2207
rect 5154 2147 5298 2163
rect 5154 2143 5264 2147
rect 5154 2109 5231 2143
rect 5398 2133 5436 2167
rect 5364 2132 5470 2133
rect 5513 2147 5570 2163
rect 5265 2109 5298 2113
rect 5154 2097 5298 2109
rect 5513 2113 5520 2147
rect 5554 2113 5570 2147
rect 5726 2133 5764 2167
rect 5798 2147 5810 2163
rect 30 2030 33 2045
rect 30 1995 67 2030
rect 30 1991 33 1995
rect 64 1957 67 1961
rect 33 1945 67 1957
rect 793 2011 827 2053
rect 793 1935 827 1977
rect 5513 1975 5570 2113
rect 5776 2097 5810 2113
rect 14004 2111 14020 2145
rect 14069 2111 14088 2145
rect 14122 2111 14154 2145
rect 14190 2111 14206 2145
rect 14256 2088 14309 2100
rect 14256 2084 14266 2088
rect 14300 2054 14309 2088
rect 14290 2050 14309 2054
rect 14256 2016 14309 2050
rect 14256 1989 14266 2016
rect 14004 1955 14020 1989
rect 14069 1955 14088 1989
rect 14122 1955 14154 1989
rect 14190 1955 14206 1989
rect 14300 1982 14309 2016
rect 14290 1955 14309 1982
rect 177 1900 193 1934
rect 227 1900 261 1934
rect 295 1900 329 1934
rect 363 1900 397 1934
rect 431 1900 465 1934
rect 499 1900 531 1934
rect 567 1900 601 1934
rect 637 1900 669 1934
rect 703 1900 719 1934
rect 33 1877 67 1889
rect 33 1803 67 1839
rect 793 1859 827 1901
rect 14256 1894 14309 1955
rect 14290 1860 14309 1894
rect 14256 1843 14309 1860
rect 14362 1843 14432 2100
rect 793 1783 827 1825
rect 14004 1799 14020 1833
rect 14069 1799 14088 1833
rect 14122 1799 14154 1833
rect 14190 1799 14206 1833
rect 33 1734 67 1754
rect 177 1744 193 1778
rect 227 1744 261 1778
rect 295 1744 329 1778
rect 363 1744 371 1778
rect 431 1744 443 1778
rect 499 1744 533 1778
rect 567 1744 601 1778
rect 635 1744 669 1778
rect 703 1744 719 1778
rect 793 1714 827 1749
rect 33 1665 67 1666
rect 33 1612 67 1631
rect 789 1707 827 1714
rect 789 1690 793 1707
rect 823 1656 827 1673
rect 789 1631 827 1656
rect 177 1588 193 1622
rect 227 1588 261 1622
rect 295 1588 329 1622
rect 363 1588 397 1622
rect 431 1588 465 1622
rect 499 1588 531 1622
rect 567 1588 601 1622
rect 637 1588 669 1622
rect 703 1588 719 1622
rect 789 1597 793 1631
rect 789 1591 827 1597
rect 33 1527 67 1562
rect 33 1477 67 1490
rect 823 1557 827 1591
rect 789 1555 827 1557
rect 789 1521 793 1555
rect 789 1491 827 1521
rect 823 1479 827 1491
rect 177 1432 193 1466
rect 227 1432 261 1466
rect 295 1432 329 1466
rect 363 1432 371 1466
rect 431 1432 443 1466
rect 499 1432 533 1466
rect 567 1432 601 1466
rect 635 1432 669 1466
rect 703 1432 719 1466
rect 789 1445 793 1457
rect 789 1433 823 1445
<< viali >>
rect 531 2648 533 2682
rect 533 2648 565 2682
rect 673 2648 703 2682
rect 703 2648 707 2682
rect 793 2654 827 2688
rect -37 2608 -3 2642
rect -37 2532 -3 2566
rect 977 2635 1011 2669
rect 1049 2635 1079 2669
rect 1079 2635 1083 2669
rect 1143 2645 1177 2649
rect 793 2579 827 2613
rect 531 2492 533 2526
rect 533 2492 565 2526
rect 603 2492 635 2526
rect 635 2492 637 2526
rect 793 2504 827 2538
rect 1143 2615 1177 2645
rect 1143 2540 1177 2570
rect 1143 2536 1177 2540
rect 869 2479 903 2513
rect 941 2479 943 2513
rect 943 2479 975 2513
rect 793 2429 827 2463
rect 288 2368 295 2402
rect 295 2368 322 2402
rect 360 2368 363 2402
rect 363 2368 394 2402
rect 30 2341 64 2345
rect 30 2311 33 2341
rect 33 2311 64 2341
rect 30 2237 33 2256
rect 33 2237 64 2256
rect 793 2354 827 2388
rect 1143 2452 1177 2456
rect 1143 2422 1177 2452
rect 977 2323 1011 2357
rect 1049 2323 1079 2357
rect 1079 2323 1083 2357
rect 1143 2347 1177 2377
rect 1143 2343 1177 2347
rect 793 2279 827 2313
rect 30 2222 64 2237
rect 531 2212 533 2246
rect 533 2212 565 2246
rect 603 2212 635 2246
rect 635 2212 637 2246
rect 30 2133 64 2167
rect 793 2204 827 2238
rect 793 2129 827 2163
rect 30 2064 64 2079
rect 30 2045 33 2064
rect 33 2045 64 2064
rect 288 2056 295 2090
rect 295 2056 322 2090
rect 360 2056 363 2090
rect 363 2056 394 2090
rect 5231 2211 5265 2245
rect 5578 2241 5612 2248
rect 5578 2214 5581 2241
rect 5581 2214 5612 2241
rect 5680 2214 5714 2248
rect 5231 2113 5264 2143
rect 5264 2113 5265 2143
rect 5364 2133 5398 2167
rect 5436 2133 5470 2167
rect 5231 2109 5265 2113
rect 5692 2133 5726 2167
rect 5764 2147 5798 2167
rect 5764 2133 5776 2147
rect 5776 2133 5798 2147
rect 30 1961 33 1991
rect 33 1961 64 1991
rect 30 1957 64 1961
rect 793 2053 827 2087
rect 793 1977 827 2011
rect 14035 2111 14054 2145
rect 14054 2111 14069 2145
rect 14154 2111 14156 2145
rect 14156 2111 14188 2145
rect 14266 2084 14300 2088
rect 14266 2054 14290 2084
rect 14290 2054 14300 2084
rect 14266 1989 14300 2016
rect 14035 1955 14054 1989
rect 14054 1955 14069 1989
rect 14154 1955 14156 1989
rect 14156 1955 14188 1989
rect 14266 1982 14290 1989
rect 14290 1982 14300 1989
rect 531 1900 533 1934
rect 533 1900 565 1934
rect 603 1900 635 1934
rect 635 1900 637 1934
rect 793 1901 827 1935
rect 33 1873 67 1877
rect 33 1843 67 1873
rect 33 1769 67 1788
rect 793 1825 827 1859
rect 14035 1799 14054 1833
rect 14054 1799 14069 1833
rect 14154 1799 14156 1833
rect 14156 1799 14188 1833
rect 33 1754 67 1769
rect 371 1744 397 1778
rect 397 1744 405 1778
rect 443 1744 465 1778
rect 465 1744 477 1778
rect 793 1749 827 1783
rect 33 1666 67 1700
rect 793 1690 827 1707
rect 793 1673 823 1690
rect 823 1673 827 1690
rect 33 1596 67 1612
rect 33 1578 67 1596
rect 531 1588 533 1622
rect 533 1588 565 1622
rect 603 1588 635 1622
rect 635 1588 637 1622
rect 793 1597 827 1631
rect 33 1493 67 1524
rect 33 1490 67 1493
rect 793 1521 827 1555
rect 371 1432 397 1466
rect 397 1432 405 1466
rect 443 1432 465 1466
rect 465 1432 477 1466
rect 793 1457 823 1479
rect 823 1457 827 1479
rect 793 1445 827 1457
<< metal1 >>
rect 34 3090 78 3122
rect -43 2642 3 2654
rect -43 2608 -37 2642
rect -3 2608 3 2642
rect -43 2566 3 2608
rect -43 2532 -37 2566
rect -3 2532 3 2566
rect -43 2520 3 2532
rect 34 2357 66 3090
rect 24 2345 70 2357
rect 24 2311 30 2345
rect 64 2311 70 2345
rect 24 2256 70 2311
rect 24 2222 30 2256
rect 64 2222 70 2256
rect 24 2167 70 2222
rect 24 2133 30 2167
rect 64 2133 70 2167
rect 24 2079 70 2133
rect 24 2045 30 2079
rect 64 2045 70 2079
rect 24 1991 70 2045
rect 24 1957 30 1991
rect 64 1957 70 1991
rect 24 1945 70 1957
tri 84 1900 98 1914 se
rect 98 1900 126 3038
rect 7935 2932 15049 2960
rect 965 2814 971 2866
rect 1023 2814 1039 2866
rect 1091 2814 1097 2866
tri 766 2688 778 2700 se
rect 778 2688 833 2700
rect 519 2682 793 2688
rect 519 2648 531 2682
rect 565 2648 673 2682
rect 707 2654 793 2682
rect 827 2654 833 2688
rect 707 2648 833 2654
rect 519 2642 833 2648
tri 758 2635 765 2642 ne
rect 765 2635 833 2642
tri 765 2615 785 2635 ne
rect 785 2615 833 2635
rect 965 2675 1096 2814
rect 965 2669 1095 2675
rect 965 2635 977 2669
rect 1011 2635 1049 2669
rect 1083 2635 1095 2669
rect 965 2629 1095 2635
rect 1137 2649 1183 2661
tri 785 2613 787 2615 ne
rect 787 2613 833 2615
rect 787 2579 793 2613
rect 827 2579 833 2613
rect 1137 2615 1143 2649
rect 1177 2615 1183 2649
rect 787 2538 833 2579
tri 1116 2570 1137 2591 se
rect 1137 2570 1183 2615
tri 1101 2555 1116 2570 se
rect 1116 2555 1143 2570
tri 1089 2543 1101 2555 se
rect 1101 2543 1143 2555
rect 519 2526 649 2532
rect 519 2492 531 2526
rect 565 2492 603 2526
rect 637 2492 649 2526
rect 276 2402 406 2408
rect 276 2368 288 2402
rect 322 2368 360 2402
rect 394 2368 406 2402
rect 276 2218 406 2368
rect 519 2246 649 2492
tri 406 2218 413 2225 sw
rect 276 2166 282 2218
rect 334 2166 355 2218
rect 407 2166 413 2218
rect 276 2163 410 2166
tri 410 2163 413 2166 nw
rect 519 2212 531 2246
rect 565 2212 603 2246
rect 637 2212 649 2246
rect 276 2090 406 2163
tri 406 2159 410 2163 nw
rect 276 2056 288 2090
rect 322 2056 360 2090
rect 394 2056 406 2090
rect 276 2050 406 2056
rect 436 2131 489 2137
rect 488 2079 489 2131
rect 436 2058 489 2079
tri 73 1889 84 1900 se
rect 84 1889 126 1900
rect 27 1881 126 1889
rect 27 1877 104 1881
rect 27 1843 33 1877
rect 67 1859 104 1877
tri 104 1859 126 1881 nw
rect 488 2006 489 2058
rect 67 1843 73 1859
rect 27 1788 73 1843
tri 73 1828 104 1859 nw
tri 431 1828 436 1833 se
rect 436 1828 489 2006
tri 428 1825 431 1828 se
rect 431 1825 489 1828
tri 409 1806 428 1825 se
rect 428 1806 489 1825
tri 402 1799 409 1806 se
rect 409 1799 489 1806
rect 27 1754 33 1788
rect 67 1754 73 1788
tri 390 1787 402 1799 se
rect 402 1787 489 1799
rect 27 1700 73 1754
rect 27 1666 33 1700
rect 67 1666 73 1700
rect 27 1612 73 1666
rect 27 1578 33 1612
rect 67 1578 73 1612
rect 27 1524 73 1578
rect 27 1490 33 1524
rect 67 1490 73 1524
rect 27 1478 73 1490
rect 359 1778 489 1787
rect 359 1744 371 1778
rect 405 1744 443 1778
rect 477 1744 489 1778
rect 359 1466 489 1744
rect 519 1934 649 2212
rect 519 1900 531 1934
rect 565 1900 603 1934
rect 637 1900 649 1934
rect 519 1622 649 1900
rect 519 1588 531 1622
rect 565 1588 603 1622
rect 637 1588 649 1622
rect 519 1582 649 1588
rect 787 2504 793 2538
rect 827 2536 833 2538
tri 833 2536 840 2543 sw
tri 1082 2536 1089 2543 se
rect 1089 2536 1143 2543
rect 1177 2536 1183 2570
rect 827 2532 840 2536
tri 840 2532 844 2536 sw
tri 1078 2532 1082 2536 se
rect 1082 2532 1183 2536
rect 827 2524 844 2532
tri 844 2524 852 2532 sw
tri 1070 2524 1078 2532 se
rect 1078 2524 1183 2532
rect 827 2519 852 2524
tri 852 2519 857 2524 sw
tri 1065 2519 1070 2524 se
rect 1070 2519 1101 2524
rect 827 2513 987 2519
rect 827 2504 869 2513
rect 787 2479 869 2504
rect 903 2479 941 2513
rect 975 2479 987 2513
rect 787 2473 987 2479
tri 1055 2509 1065 2519 se
rect 1065 2509 1101 2519
rect 787 2463 839 2473
rect 787 2429 793 2463
rect 827 2456 839 2463
tri 839 2456 856 2473 nw
rect 827 2429 833 2456
tri 833 2450 839 2456 nw
rect 787 2388 833 2429
rect 787 2354 793 2388
rect 827 2354 833 2388
tri 1043 2377 1055 2389 se
rect 1055 2377 1101 2509
tri 1101 2488 1137 2524 nw
tri 1029 2363 1043 2377 se
rect 1043 2363 1101 2377
tri 923 2357 929 2363 se
rect 929 2357 1101 2363
rect 787 2313 833 2354
tri 889 2323 923 2357 se
rect 923 2323 977 2357
rect 1011 2323 1049 2357
rect 1083 2323 1101 2357
rect 1137 2456 1183 2468
rect 1137 2422 1143 2456
rect 1177 2422 1183 2456
rect 1137 2377 1183 2422
rect 1137 2343 1143 2377
rect 1177 2343 1183 2377
rect 1137 2331 1183 2343
rect 787 2279 793 2313
rect 827 2279 833 2313
rect 787 2238 833 2279
rect 787 2204 793 2238
rect 827 2204 833 2238
rect 787 2163 833 2204
tri 886 2320 889 2323 se
rect 889 2320 1101 2323
rect 886 2317 1101 2320
rect 886 2305 953 2317
tri 953 2305 965 2317 nw
rect 886 2299 938 2305
tri 938 2290 953 2305 nw
rect 886 2226 938 2247
rect 5154 2205 5160 2257
rect 5212 2205 5224 2257
rect 5276 2205 5282 2257
rect 5565 2205 5571 2257
rect 5623 2205 5639 2257
rect 5691 2248 5707 2257
rect 5691 2205 5707 2214
rect 5759 2205 5765 2257
rect 886 2168 938 2174
rect 787 2129 793 2163
rect 827 2129 833 2163
rect 787 2087 833 2129
rect 5225 2143 5271 2205
rect 5225 2109 5231 2143
rect 5265 2109 5271 2143
rect 5352 2123 5358 2175
rect 5410 2123 5422 2175
rect 5474 2173 5480 2175
rect 5474 2127 5482 2173
rect 5474 2123 5480 2127
rect 5680 2123 5686 2175
rect 5738 2123 5750 2175
rect 5802 2173 5808 2175
rect 5802 2127 5810 2173
rect 5802 2123 5808 2127
rect 5225 2097 5271 2109
rect 7935 2095 7963 2932
rect 14256 2448 14980 2477
rect 8012 2247 8064 2253
rect 8012 2183 8064 2195
tri 13955 2145 13961 2151 se
rect 13961 2145 14200 2151
rect 8012 2125 8064 2131
tri 13935 2125 13955 2145 se
rect 13955 2125 14035 2145
tri 13926 2116 13935 2125 se
rect 13935 2116 14035 2125
rect 13926 2111 14035 2116
rect 14069 2111 14154 2145
rect 14188 2111 14200 2145
rect 13926 2105 14200 2111
rect 13926 2095 14038 2105
tri 14038 2095 14048 2105 nw
rect 787 2053 793 2087
rect 827 2053 833 2087
rect 787 2011 833 2053
rect 787 1977 793 2011
rect 827 1977 833 2011
rect 787 1935 833 1977
rect 787 1901 793 1935
rect 827 1901 833 1935
rect 787 1859 833 1901
rect 787 1825 793 1859
rect 827 1825 833 1859
rect 787 1783 833 1825
rect 13926 2088 14031 2095
tri 14031 2088 14038 2095 nw
rect 14256 2088 14326 2448
rect 15021 2414 15049 2932
rect 13926 2054 13997 2088
tri 13997 2054 14031 2088 nw
rect 14256 2054 14266 2088
rect 14300 2054 14326 2088
rect 13926 1839 13991 2054
tri 13991 2048 13997 2054 nw
rect 14256 2016 14326 2054
rect 14023 1989 14200 1995
rect 14023 1955 14035 1989
rect 14069 1955 14154 1989
rect 14188 1955 14200 1989
rect 14256 1982 14266 2016
rect 14300 1982 14326 2016
rect 14256 1970 14326 1982
rect 14362 2382 15049 2414
rect 14362 1970 14432 2382
rect 14688 1993 15108 2027
rect 14023 1922 14200 1955
rect 14688 1922 14722 1993
rect 14023 1888 14722 1922
tri 13991 1839 14017 1865 sw
rect 13926 1833 14200 1839
rect 13926 1821 14035 1833
tri 13926 1799 13948 1821 ne
rect 13948 1799 14035 1821
rect 14069 1799 14154 1833
rect 14188 1799 14200 1833
tri 13948 1793 13954 1799 ne
rect 13954 1793 14200 1799
rect 787 1749 793 1783
rect 827 1749 833 1783
rect 787 1707 833 1749
rect 787 1673 793 1707
rect 827 1673 833 1707
rect 787 1631 833 1673
rect 787 1597 793 1631
rect 827 1597 833 1631
rect 359 1432 371 1466
rect 405 1432 443 1466
rect 477 1432 489 1466
rect 787 1555 833 1597
rect 787 1521 793 1555
rect 827 1521 833 1555
rect 787 1479 833 1521
rect 787 1445 793 1479
rect 827 1445 833 1479
rect 787 1433 833 1445
rect 359 1426 489 1432
<< via1 >>
rect 971 2814 1023 2866
rect 1039 2814 1091 2866
rect 282 2166 334 2218
rect 355 2166 407 2218
rect 436 2079 488 2131
rect 436 2006 488 2058
rect 886 2247 938 2299
rect 886 2174 938 2226
rect 5160 2205 5212 2257
rect 5224 2245 5276 2257
rect 5224 2211 5231 2245
rect 5231 2211 5265 2245
rect 5265 2211 5276 2245
rect 5224 2205 5276 2211
rect 5571 2248 5623 2257
rect 5571 2214 5578 2248
rect 5578 2214 5612 2248
rect 5612 2214 5623 2248
rect 5571 2205 5623 2214
rect 5639 2248 5691 2257
rect 5707 2248 5759 2257
rect 5639 2214 5680 2248
rect 5680 2214 5691 2248
rect 5707 2214 5714 2248
rect 5714 2214 5759 2248
rect 5639 2205 5691 2214
rect 5707 2205 5759 2214
rect 5358 2167 5410 2175
rect 5358 2133 5364 2167
rect 5364 2133 5398 2167
rect 5398 2133 5410 2167
rect 5358 2123 5410 2133
rect 5422 2167 5474 2175
rect 5422 2133 5436 2167
rect 5436 2133 5470 2167
rect 5470 2133 5474 2167
rect 5422 2123 5474 2133
rect 5686 2167 5738 2175
rect 5686 2133 5692 2167
rect 5692 2133 5726 2167
rect 5726 2133 5738 2167
rect 5686 2123 5738 2133
rect 5750 2167 5802 2175
rect 5750 2133 5764 2167
rect 5764 2133 5798 2167
rect 5798 2133 5802 2167
rect 5750 2123 5802 2133
rect 8012 2195 8064 2247
rect 8012 2131 8064 2183
<< metal2 >>
rect 965 2814 971 2866
rect 1023 2814 1039 2866
rect 1091 2836 7720 2866
rect 1091 2814 1097 2836
rect 886 2299 938 2305
rect 886 2226 938 2247
tri 1109 2232 1134 2257 se
rect 1134 2232 5160 2257
rect 276 2166 282 2218
rect 334 2166 355 2218
rect 407 2174 886 2218
tri 1095 2218 1109 2232 se
rect 1109 2218 5160 2232
rect 938 2205 5160 2218
rect 5212 2205 5224 2257
rect 5276 2205 5571 2257
rect 5623 2205 5639 2257
rect 5691 2205 5707 2257
rect 5759 2247 6377 2257
tri 6377 2247 6387 2257 sw
rect 8012 2247 8064 2253
rect 5759 2232 6387 2247
tri 6387 2232 6402 2247 sw
rect 5759 2205 6402 2232
rect 938 2195 1163 2205
tri 1163 2195 1173 2205 nw
tri 6364 2195 6374 2205 ne
rect 6374 2195 6402 2205
tri 6402 2195 6439 2232 sw
rect 938 2183 1151 2195
tri 1151 2183 1163 2195 nw
tri 6374 2183 6386 2195 ne
rect 6386 2183 6439 2195
tri 6439 2183 6451 2195 sw
tri 7152 2183 7162 2193 se
rect 7162 2183 7559 2193
tri 7559 2183 7569 2193 sw
rect 8012 2183 8064 2195
rect 938 2175 1143 2183
tri 1143 2175 1151 2183 nw
tri 6386 2175 6394 2183 ne
rect 6394 2175 6451 2183
rect 938 2174 1135 2175
rect 407 2167 1135 2174
tri 1135 2167 1143 2175 nw
tri 1280 2167 1288 2175 se
rect 1288 2167 5358 2175
rect 407 2166 1134 2167
tri 1134 2166 1135 2167 nw
tri 1279 2166 1280 2167 se
rect 1280 2166 5358 2167
tri 1250 2137 1279 2166 se
rect 1279 2137 5358 2166
rect 436 2131 5358 2137
rect 488 2123 5358 2131
rect 5410 2123 5422 2175
rect 5474 2123 5686 2175
rect 5738 2123 5750 2175
rect 5802 2123 5810 2175
tri 6394 2167 6402 2175 ne
rect 6402 2167 6451 2175
tri 6451 2167 6467 2183 sw
tri 7136 2167 7152 2183 se
rect 7152 2167 7569 2183
tri 7569 2167 7585 2183 sw
tri 6402 2166 6403 2167 ne
rect 6403 2166 7585 2167
tri 6403 2131 6438 2166 ne
rect 6438 2158 7585 2166
tri 7585 2158 7594 2167 sw
rect 6438 2155 8012 2158
rect 6438 2131 7176 2155
tri 7176 2131 7200 2155 nw
tri 7536 2131 7560 2155 ne
rect 7560 2131 8012 2155
tri 6438 2123 6446 2131 ne
rect 6446 2125 7170 2131
tri 7170 2125 7176 2131 nw
tri 7560 2125 7566 2131 ne
rect 7566 2125 8064 2131
rect 6446 2123 7167 2125
rect 488 2122 1326 2123
tri 1326 2122 1327 2123 nw
tri 6446 2122 6447 2123 ne
rect 6447 2122 7167 2123
tri 7167 2122 7170 2125 nw
rect 488 2085 1289 2122
tri 1289 2085 1326 2122 nw
rect 436 2058 488 2079
rect 436 2000 488 2006
use sky130_fd_pr__nfet_01v8__example_55959141808483  sky130_fd_pr__nfet_01v8__example_55959141808483_0
timestamp 1663361622
transform 0 -1 715 -1 0 2357
box -1 0 881 1
use sky130_fd_pr__nfet_01v8__example_55959141808484  sky130_fd_pr__nfet_01v8__example_55959141808484_0
timestamp 1663361622
transform 0 -1 715 -1 0 2637
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808485  sky130_fd_pr__nfet_01v8__example_55959141808485_0
timestamp 1663361622
transform 0 1 897 1 0 2368
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808482  sky130_fd_pr__pfet_01v8__example_55959141808482_0
timestamp 1663361622
transform -1 0 5765 0 -1 2159
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808482  sky130_fd_pr__pfet_01v8__example_55959141808482_1
timestamp 1663361622
transform -1 0 5509 0 -1 2159
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808512  sky130_fd_pr__pfet_01v8__example_55959141808512_0
timestamp 1663361622
transform 0 1 14008 -1 0 2100
box -1 0 257 1
<< labels >>
flabel comment s 57 2394 57 2394 0 FreeSans 280 90 0 0 IN_B
flabel comment s 115 2434 115 2434 0 FreeSans 280 90 0 0 IN
<< properties >>
string GDS_END 29588372
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 29571158
<< end >>
