magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 1 5 1 5 6 DRAIN
port 2 nsew
rlabel  s 0 5 1 6 4 GATE
port 3 nsew
rlabel  s 1 0 1 5 6 SOURCE
port 4 nsew
rlabel  s 0 0 0 5 4 SOURCE
port 4 nsew
rlabel  s 0 0 1 0 2 SOURCE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 1 6
string LEFview TRUE
<< end >>
