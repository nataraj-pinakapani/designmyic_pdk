magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 160 1251
rect 560 403 867 865
rect 1267 493 2274 1251
rect 1960 377 2274 493
<< pwell >>
rect -26 1585 2234 1671
rect 637 1195 1051 1585
rect 1781 1345 2204 1585
rect 1018 345 1900 433
rect 571 43 1900 345
rect -26 -43 2234 43
<< scnmos >>
rect 656 151 686 319
rect 742 151 772 319
<< scpmoshvt >>
rect 656 439 686 607
rect 742 439 772 607
<< mvnmos >>
rect 716 1221 816 1521
rect 872 1221 972 1521
rect 1860 1371 1960 1521
rect 2025 1371 2125 1521
rect 1097 107 1197 407
rect 1253 107 1353 407
rect 1565 107 1665 407
rect 1721 107 1821 407
<< mvpmos >>
rect 1400 885 1500 1185
rect 1565 885 1665 1185
rect 1860 885 1960 1185
rect 2025 885 2125 1185
rect 1406 563 1606 647
rect 1694 563 1894 647
rect 1982 563 2082 647
<< ndiff >>
rect 597 299 656 319
rect 597 265 611 299
rect 645 265 656 299
rect 597 197 656 265
rect 597 163 611 197
rect 645 163 656 197
rect 597 151 656 163
rect 686 299 742 319
rect 686 265 697 299
rect 731 265 742 299
rect 686 193 742 265
rect 686 159 697 193
rect 731 159 742 193
rect 686 151 742 159
rect 772 299 831 319
rect 772 265 783 299
rect 817 265 831 299
rect 772 197 831 265
rect 772 163 783 197
rect 817 163 831 197
rect 772 151 831 163
<< pdiff >>
rect 597 595 656 607
rect 597 561 611 595
rect 645 561 656 595
rect 597 483 656 561
rect 597 449 611 483
rect 645 449 656 483
rect 597 439 656 449
rect 686 595 742 607
rect 686 561 697 595
rect 731 561 742 595
rect 686 483 742 561
rect 686 449 697 483
rect 731 449 742 483
rect 686 439 742 449
rect 772 565 831 607
rect 772 531 783 565
rect 817 531 831 565
rect 772 483 831 531
rect 772 449 783 483
rect 817 449 831 483
rect 772 439 831 449
<< mvndiff >>
rect 663 1509 716 1521
rect 663 1475 671 1509
rect 705 1475 716 1509
rect 663 1429 716 1475
rect 663 1395 671 1429
rect 705 1395 716 1429
rect 663 1347 716 1395
rect 663 1313 671 1347
rect 705 1313 716 1347
rect 663 1267 716 1313
rect 663 1233 671 1267
rect 705 1233 716 1267
rect 663 1221 716 1233
rect 816 1509 872 1521
rect 816 1475 827 1509
rect 861 1475 872 1509
rect 816 1429 872 1475
rect 816 1395 827 1429
rect 861 1395 872 1429
rect 816 1347 872 1395
rect 816 1313 827 1347
rect 861 1313 872 1347
rect 816 1267 872 1313
rect 816 1233 827 1267
rect 861 1233 872 1267
rect 816 1221 872 1233
rect 972 1509 1025 1521
rect 972 1475 983 1509
rect 1017 1475 1025 1509
rect 972 1429 1025 1475
rect 972 1395 983 1429
rect 1017 1395 1025 1429
rect 972 1347 1025 1395
rect 1807 1509 1860 1521
rect 1807 1475 1815 1509
rect 1849 1475 1860 1509
rect 1807 1417 1860 1475
rect 972 1313 983 1347
rect 1017 1313 1025 1347
rect 972 1267 1025 1313
rect 1807 1383 1815 1417
rect 1849 1383 1860 1417
rect 1807 1371 1860 1383
rect 1960 1509 2025 1521
rect 1960 1475 1980 1509
rect 2014 1475 2025 1509
rect 1960 1417 2025 1475
rect 1960 1383 1980 1417
rect 2014 1383 2025 1417
rect 1960 1371 2025 1383
rect 2125 1509 2178 1521
rect 2125 1475 2136 1509
rect 2170 1475 2178 1509
rect 2125 1417 2178 1475
rect 2125 1383 2136 1417
rect 2170 1383 2178 1417
rect 2125 1371 2178 1383
rect 972 1233 983 1267
rect 1017 1233 1025 1267
rect 972 1221 1025 1233
rect 1044 395 1097 407
rect 1044 361 1052 395
rect 1086 361 1097 395
rect 1044 315 1097 361
rect 1044 281 1052 315
rect 1086 281 1097 315
rect 1044 233 1097 281
rect 1044 199 1052 233
rect 1086 199 1097 233
rect 1044 153 1097 199
rect 1044 119 1052 153
rect 1086 119 1097 153
rect 1044 107 1097 119
rect 1197 395 1253 407
rect 1197 361 1208 395
rect 1242 361 1253 395
rect 1197 315 1253 361
rect 1197 281 1208 315
rect 1242 281 1253 315
rect 1197 233 1253 281
rect 1197 199 1208 233
rect 1242 199 1253 233
rect 1197 153 1253 199
rect 1197 119 1208 153
rect 1242 119 1253 153
rect 1197 107 1253 119
rect 1353 395 1406 407
rect 1353 361 1364 395
rect 1398 361 1406 395
rect 1353 315 1406 361
rect 1353 281 1364 315
rect 1398 281 1406 315
rect 1353 233 1406 281
rect 1353 199 1364 233
rect 1398 199 1406 233
rect 1353 153 1406 199
rect 1353 119 1364 153
rect 1398 119 1406 153
rect 1353 107 1406 119
rect 1512 395 1565 407
rect 1512 361 1520 395
rect 1554 361 1565 395
rect 1512 315 1565 361
rect 1512 281 1520 315
rect 1554 281 1565 315
rect 1512 233 1565 281
rect 1512 199 1520 233
rect 1554 199 1565 233
rect 1512 153 1565 199
rect 1512 119 1520 153
rect 1554 119 1565 153
rect 1512 107 1565 119
rect 1665 395 1721 407
rect 1665 361 1676 395
rect 1710 361 1721 395
rect 1665 315 1721 361
rect 1665 281 1676 315
rect 1710 281 1721 315
rect 1665 233 1721 281
rect 1665 199 1676 233
rect 1710 199 1721 233
rect 1665 153 1721 199
rect 1665 119 1676 153
rect 1710 119 1721 153
rect 1665 107 1721 119
rect 1821 395 1874 407
rect 1821 361 1832 395
rect 1866 361 1874 395
rect 1821 315 1874 361
rect 1821 281 1832 315
rect 1866 281 1874 315
rect 1821 233 1874 281
rect 1821 199 1832 233
rect 1866 199 1874 233
rect 1821 153 1874 199
rect 1821 119 1832 153
rect 1866 119 1874 153
rect 1821 107 1874 119
<< mvpdiff >>
rect 1347 1173 1400 1185
rect 1347 1139 1355 1173
rect 1389 1139 1400 1173
rect 1347 1093 1400 1139
rect 1347 1059 1355 1093
rect 1389 1059 1400 1093
rect 1347 1011 1400 1059
rect 1347 977 1355 1011
rect 1389 977 1400 1011
rect 1347 931 1400 977
rect 1347 897 1355 931
rect 1389 897 1400 931
rect 1347 885 1400 897
rect 1500 1173 1565 1185
rect 1500 1139 1520 1173
rect 1554 1139 1565 1173
rect 1500 1093 1565 1139
rect 1500 1059 1520 1093
rect 1554 1059 1565 1093
rect 1500 1011 1565 1059
rect 1500 977 1520 1011
rect 1554 977 1565 1011
rect 1500 931 1565 977
rect 1500 897 1520 931
rect 1554 897 1565 931
rect 1500 885 1565 897
rect 1665 1173 1718 1185
rect 1665 1139 1676 1173
rect 1710 1139 1718 1173
rect 1665 1093 1718 1139
rect 1665 1059 1676 1093
rect 1710 1059 1718 1093
rect 1665 1011 1718 1059
rect 1665 977 1676 1011
rect 1710 977 1718 1011
rect 1665 931 1718 977
rect 1665 897 1676 931
rect 1710 897 1718 931
rect 1665 885 1718 897
rect 1807 1173 1860 1185
rect 1807 1139 1815 1173
rect 1849 1139 1860 1173
rect 1807 1093 1860 1139
rect 1807 1059 1815 1093
rect 1849 1059 1860 1093
rect 1807 1011 1860 1059
rect 1807 977 1815 1011
rect 1849 977 1860 1011
rect 1807 931 1860 977
rect 1807 897 1815 931
rect 1849 897 1860 931
rect 1807 885 1860 897
rect 1960 1173 2025 1185
rect 1960 1139 1980 1173
rect 2014 1139 2025 1173
rect 1960 1093 2025 1139
rect 1960 1059 1980 1093
rect 2014 1059 2025 1093
rect 1960 1011 2025 1059
rect 1960 977 1980 1011
rect 2014 977 2025 1011
rect 1960 931 2025 977
rect 1960 897 1980 931
rect 2014 897 2025 931
rect 1960 885 2025 897
rect 2125 1173 2178 1185
rect 2125 1139 2136 1173
rect 2170 1139 2178 1173
rect 2125 1093 2178 1139
rect 2125 1059 2136 1093
rect 2170 1059 2178 1093
rect 2125 1011 2178 1059
rect 2125 977 2136 1011
rect 2170 977 2178 1011
rect 2125 931 2178 977
rect 2125 897 2136 931
rect 2170 897 2178 931
rect 2125 885 2178 897
rect 1333 677 1391 689
rect 1333 643 1345 677
rect 1379 647 1391 677
rect 1621 677 1679 689
rect 1621 647 1633 677
rect 1379 643 1406 647
rect 1333 609 1406 643
rect 1333 575 1345 609
rect 1379 575 1406 609
rect 1333 563 1406 575
rect 1606 643 1633 647
rect 1667 647 1679 677
rect 1909 677 1967 689
rect 1909 647 1921 677
rect 1667 643 1694 647
rect 1606 609 1694 643
rect 1606 575 1633 609
rect 1667 575 1694 609
rect 1606 563 1694 575
rect 1894 643 1921 647
rect 1955 647 1967 677
rect 2097 677 2155 689
rect 2097 647 2109 677
rect 1955 643 1982 647
rect 1894 609 1982 643
rect 1894 575 1921 609
rect 1955 575 1982 609
rect 1894 563 1982 575
rect 2082 643 2109 647
rect 2143 643 2155 677
rect 2082 609 2155 643
rect 2082 575 2109 609
rect 2143 575 2155 609
rect 2082 563 2155 575
<< ndiffc >>
rect 611 265 645 299
rect 611 163 645 197
rect 697 265 731 299
rect 697 159 731 193
rect 783 265 817 299
rect 783 163 817 197
<< pdiffc >>
rect 611 561 645 595
rect 611 449 645 483
rect 697 561 731 595
rect 697 449 731 483
rect 783 531 817 565
rect 783 449 817 483
<< mvndiffc >>
rect 671 1475 705 1509
rect 671 1395 705 1429
rect 671 1313 705 1347
rect 671 1233 705 1267
rect 827 1475 861 1509
rect 827 1395 861 1429
rect 827 1313 861 1347
rect 827 1233 861 1267
rect 983 1475 1017 1509
rect 983 1395 1017 1429
rect 1815 1475 1849 1509
rect 983 1313 1017 1347
rect 1815 1383 1849 1417
rect 1980 1475 2014 1509
rect 1980 1383 2014 1417
rect 2136 1475 2170 1509
rect 2136 1383 2170 1417
rect 983 1233 1017 1267
rect 1052 361 1086 395
rect 1052 281 1086 315
rect 1052 199 1086 233
rect 1052 119 1086 153
rect 1208 361 1242 395
rect 1208 281 1242 315
rect 1208 199 1242 233
rect 1208 119 1242 153
rect 1364 361 1398 395
rect 1364 281 1398 315
rect 1364 199 1398 233
rect 1364 119 1398 153
rect 1520 361 1554 395
rect 1520 281 1554 315
rect 1520 199 1554 233
rect 1520 119 1554 153
rect 1676 361 1710 395
rect 1676 281 1710 315
rect 1676 199 1710 233
rect 1676 119 1710 153
rect 1832 361 1866 395
rect 1832 281 1866 315
rect 1832 199 1866 233
rect 1832 119 1866 153
<< mvpdiffc >>
rect 1355 1139 1389 1173
rect 1355 1059 1389 1093
rect 1355 977 1389 1011
rect 1355 897 1389 931
rect 1520 1139 1554 1173
rect 1520 1059 1554 1093
rect 1520 977 1554 1011
rect 1520 897 1554 931
rect 1676 1139 1710 1173
rect 1676 1059 1710 1093
rect 1676 977 1710 1011
rect 1676 897 1710 931
rect 1815 1139 1849 1173
rect 1815 1059 1849 1093
rect 1815 977 1849 1011
rect 1815 897 1849 931
rect 1980 1139 2014 1173
rect 1980 1059 2014 1093
rect 1980 977 2014 1011
rect 1980 897 2014 931
rect 2136 1139 2170 1173
rect 2136 1059 2170 1093
rect 2136 977 2170 1011
rect 2136 897 2170 931
rect 1345 643 1379 677
rect 1345 575 1379 609
rect 1633 643 1667 677
rect 1633 575 1667 609
rect 1921 643 1955 677
rect 1921 575 1955 609
rect 2109 643 2143 677
rect 2109 575 2143 609
<< nsubdiff >>
rect 653 824 831 829
rect 653 790 677 824
rect 711 790 773 824
rect 807 790 831 824
rect 653 714 831 790
rect 653 680 677 714
rect 711 680 773 714
rect 807 680 831 714
rect 653 661 831 680
<< mvpsubdiff >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2208 1645
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 94 831
rect 1639 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1849 831
rect 2112 797 2143 831
rect 2177 797 2208 831
<< nsubdiffcont >>
rect 677 790 711 824
rect 773 790 807 824
rect 677 680 711 714
rect 773 680 807 714
<< mvpsubdiffcont >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 2143 797 2177 831
<< poly >>
rect 716 1521 816 1547
rect 872 1521 972 1547
rect 1860 1521 1960 1547
rect 2025 1521 2125 1547
rect 1707 1375 1773 1391
rect 1707 1341 1723 1375
rect 1757 1341 1773 1375
rect 1707 1323 1773 1341
rect 1860 1345 1960 1371
rect 1860 1323 1944 1345
rect 1707 1307 1944 1323
rect 2025 1311 2125 1371
rect 716 1199 816 1221
rect 872 1199 972 1221
rect 573 1133 972 1199
rect 1400 1211 1665 1277
rect 1707 1273 1723 1307
rect 1757 1273 1944 1307
rect 1707 1257 1944 1273
rect 1400 1185 1500 1211
rect 1565 1185 1665 1211
rect 1860 1211 1944 1257
rect 1986 1295 2125 1311
rect 1986 1261 2002 1295
rect 2036 1261 2070 1295
rect 2104 1261 2125 1295
rect 1986 1245 2125 1261
rect 1860 1185 1960 1211
rect 2025 1185 2125 1245
rect 573 1083 639 1133
rect 573 1049 589 1083
rect 623 1049 639 1083
rect 573 1015 639 1049
rect 573 981 589 1015
rect 623 981 639 1015
rect 573 947 639 981
rect 573 913 589 947
rect 623 913 639 947
rect 573 897 639 913
rect 1400 870 1500 885
rect 1565 870 1665 885
rect 1400 842 1665 870
rect 1860 857 1960 885
rect 2025 870 2125 885
rect 1400 827 1628 842
rect 1400 793 1435 827
rect 1469 793 1503 827
rect 1537 793 1628 827
rect 1400 777 1628 793
rect 1860 786 1916 857
rect 2002 842 2125 870
rect 2002 815 2101 842
rect 1694 704 1916 786
rect 1982 781 2101 815
rect 1406 647 1606 673
rect 656 607 686 633
rect 742 607 772 633
rect 499 424 565 440
rect 1694 647 1894 704
rect 1982 647 2082 781
rect 1406 495 1606 563
rect 1694 537 1894 563
rect 1982 495 2082 563
rect 956 479 1353 495
rect 956 445 972 479
rect 1006 445 1040 479
rect 1074 445 1108 479
rect 1142 445 1353 479
rect 499 390 515 424
rect 549 407 565 424
rect 656 407 686 439
rect 742 407 772 439
rect 956 429 1353 445
rect 1406 429 2082 495
rect 1097 407 1197 429
rect 1253 407 1353 429
rect 1565 407 1665 429
rect 1721 407 1821 429
rect 549 390 686 407
rect 499 356 686 390
rect 499 322 515 356
rect 549 341 686 356
rect 728 391 862 407
rect 728 357 744 391
rect 778 357 812 391
rect 846 357 862 391
rect 728 341 862 357
rect 549 322 565 341
rect 499 306 565 322
rect 656 319 686 341
rect 742 319 772 341
rect 656 125 686 151
rect 742 125 772 151
rect 1097 81 1197 107
rect 1253 81 1353 107
rect 1565 81 1665 107
rect 1721 81 1821 107
<< polycont >>
rect 1723 1341 1757 1375
rect 1723 1273 1757 1307
rect 2002 1261 2036 1295
rect 2070 1261 2104 1295
rect 589 1049 623 1083
rect 589 981 623 1015
rect 589 913 623 947
rect 1435 793 1469 827
rect 1503 793 1537 827
rect 972 445 1006 479
rect 1040 445 1074 479
rect 1108 445 1142 479
rect 515 390 549 424
rect 515 322 549 356
rect 744 357 778 391
rect 812 357 846 391
<< locali >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2208 1645
rect 629 1543 1059 1577
rect 629 1509 635 1543
rect 669 1509 707 1543
rect 741 1509 747 1543
rect 941 1509 947 1543
rect 981 1509 1019 1543
rect 1053 1509 1059 1543
rect 1938 1543 2056 1549
rect 629 1475 671 1509
rect 705 1475 747 1509
rect 629 1429 747 1475
rect 629 1395 671 1429
rect 705 1395 747 1429
rect 629 1347 747 1395
rect 629 1313 671 1347
rect 705 1313 747 1347
rect 629 1267 747 1313
rect 629 1233 671 1267
rect 705 1233 747 1267
rect 811 1475 827 1509
rect 861 1475 877 1509
rect 811 1429 877 1475
rect 811 1395 827 1429
rect 861 1395 877 1429
rect 811 1347 877 1395
rect 811 1313 827 1347
rect 861 1313 877 1347
rect 811 1267 877 1313
rect 811 1233 827 1267
rect 861 1233 877 1267
rect 941 1475 983 1509
rect 1017 1475 1059 1509
rect 941 1429 1059 1475
rect 941 1395 983 1429
rect 1017 1395 1059 1429
rect 941 1347 1059 1395
rect 1799 1509 1865 1525
rect 1799 1475 1815 1509
rect 1849 1475 1865 1509
rect 1799 1417 1865 1475
rect 941 1313 983 1347
rect 1017 1313 1059 1347
rect 1707 1375 1763 1391
rect 1707 1341 1723 1375
rect 1757 1341 1763 1375
rect 1707 1323 1763 1341
rect 941 1267 1059 1313
rect 941 1233 983 1267
rect 1017 1233 1059 1267
rect 1339 1307 1763 1323
rect 1339 1273 1723 1307
rect 1757 1273 1763 1307
rect 1339 1257 1763 1273
rect 1799 1383 1815 1417
rect 1849 1383 1865 1417
rect 1799 1311 1865 1383
rect 1938 1509 1944 1543
rect 1978 1509 2016 1543
rect 2050 1509 2056 1543
rect 1938 1475 1980 1509
rect 2014 1475 2056 1509
rect 1938 1417 2056 1475
rect 1938 1383 1980 1417
rect 2014 1383 2056 1417
rect 1938 1367 2056 1383
rect 2120 1509 2186 1525
rect 2120 1475 2136 1509
rect 2170 1475 2186 1509
rect 2120 1417 2186 1475
rect 2120 1383 2136 1417
rect 2170 1383 2186 1417
rect 2120 1345 2186 1383
rect 1799 1295 2104 1311
rect 1799 1261 2002 1295
rect 2036 1261 2070 1295
rect 811 1199 877 1233
rect 1339 1199 1405 1257
rect 811 1173 1405 1199
rect 811 1139 1355 1173
rect 1389 1139 1405 1173
rect 811 1133 1405 1139
rect 577 1083 635 1099
rect 577 1049 589 1083
rect 623 1049 635 1083
rect 577 1015 635 1049
rect 577 981 589 1015
rect 623 981 635 1015
rect 577 947 635 981
rect 1339 1093 1405 1133
rect 1339 1059 1355 1093
rect 1389 1059 1405 1093
rect 1339 1011 1405 1059
rect 1339 977 1355 1011
rect 1389 977 1405 1011
rect 1339 947 1405 977
rect 577 913 589 947
rect 623 913 635 947
rect 0 797 31 831
rect 65 797 160 831
rect 577 611 635 913
rect 1313 931 1405 947
rect 1313 897 1355 931
rect 1389 897 1405 931
rect 1313 881 1405 897
rect 1478 1173 1596 1189
rect 1478 1139 1520 1173
rect 1554 1139 1596 1173
rect 1478 1093 1596 1139
rect 1478 1059 1520 1093
rect 1554 1059 1596 1093
rect 1478 1011 1596 1059
rect 1478 977 1520 1011
rect 1554 977 1596 1011
rect 1478 933 1596 977
rect 1478 899 1484 933
rect 1518 931 1556 933
rect 1518 899 1520 931
rect 1478 897 1520 899
rect 1554 899 1556 931
rect 1590 899 1596 933
rect 1554 897 1596 899
rect 1478 881 1596 897
rect 1660 1173 1726 1257
rect 1660 1139 1676 1173
rect 1710 1139 1726 1173
rect 1660 1093 1726 1139
rect 1660 1059 1676 1093
rect 1710 1059 1726 1093
rect 1660 1011 1726 1059
rect 1660 977 1676 1011
rect 1710 977 1726 1011
rect 1660 931 1726 977
rect 1660 897 1676 931
rect 1710 897 1726 931
rect 1660 881 1726 897
rect 1799 1245 2104 1261
rect 1799 1173 1865 1245
rect 2138 1211 2186 1345
rect 1799 1139 1815 1173
rect 1849 1139 1865 1173
rect 1799 1093 1865 1139
rect 1799 1059 1815 1093
rect 1849 1059 1865 1093
rect 1799 1011 1865 1059
rect 1799 977 1815 1011
rect 1849 977 1865 1011
rect 1799 931 1865 977
rect 1799 897 1815 931
rect 1849 897 1865 931
rect 1799 881 1865 897
rect 1938 1173 2056 1189
rect 1938 1139 1980 1173
rect 2014 1139 2056 1173
rect 1938 1093 2056 1139
rect 1938 1059 1980 1093
rect 2014 1059 2056 1093
rect 1938 1011 2056 1059
rect 1938 977 1980 1011
rect 2014 977 2056 1011
rect 1938 933 2056 977
rect 1938 899 1944 933
rect 1978 931 2016 933
rect 1978 899 1980 931
rect 1938 897 1980 899
rect 2014 899 2016 931
rect 2050 899 2056 933
rect 2014 897 2056 899
rect 1938 881 2056 897
rect 2120 1173 2186 1211
rect 2120 1139 2136 1173
rect 2170 1139 2186 1173
rect 2120 1093 2186 1139
rect 2120 1059 2136 1093
rect 2170 1059 2186 1093
rect 2120 1011 2186 1059
rect 2120 977 2136 1011
rect 2170 977 2186 1011
rect 2120 931 2186 977
rect 2120 897 2136 931
rect 2170 897 2186 931
rect 2120 881 2186 897
rect 669 824 823 840
rect 669 790 677 824
rect 711 790 773 824
rect 807 790 823 824
rect 669 714 823 790
rect 669 680 677 714
rect 711 680 773 714
rect 807 680 823 714
rect 669 655 823 680
rect 669 645 769 655
rect 687 644 769 645
rect 577 595 653 611
rect 577 561 611 595
rect 645 561 653 595
rect 577 553 653 561
rect 595 483 653 553
rect 595 449 611 483
rect 645 449 653 483
rect 499 424 561 440
rect 499 390 515 424
rect 549 390 561 424
rect 499 356 561 390
rect 499 322 515 356
rect 549 322 561 356
rect 499 306 561 322
rect 595 399 653 449
rect 687 610 697 644
rect 731 621 769 644
rect 803 621 823 655
rect 731 615 823 621
rect 1313 677 1379 881
rect 1313 643 1345 677
rect 731 610 741 615
rect 687 595 741 610
rect 687 561 697 595
rect 731 561 741 595
rect 1313 609 1379 643
rect 687 483 741 561
rect 687 449 697 483
rect 731 449 741 483
rect 687 433 741 449
rect 775 565 837 581
rect 775 531 783 565
rect 817 531 837 565
rect 1313 575 1345 609
rect 1313 559 1379 575
rect 1419 827 1553 843
rect 1419 793 1435 827
rect 1469 793 1503 827
rect 1537 793 1553 827
rect 1647 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2208 831
rect 775 495 837 531
rect 1419 541 1553 793
rect 1591 729 1709 741
rect 1591 695 1597 729
rect 1631 695 1669 729
rect 1703 695 1709 729
rect 1591 677 1709 695
rect 2025 729 2143 741
rect 2025 695 2031 729
rect 2065 695 2103 729
rect 2137 695 2143 729
rect 1591 643 1633 677
rect 1667 643 1709 677
rect 1591 609 1709 643
rect 1591 575 1633 609
rect 1667 575 1709 609
rect 1783 677 1967 693
rect 1783 643 1921 677
rect 1955 643 1967 677
rect 1783 609 1967 643
rect 1783 575 1921 609
rect 1955 575 1967 609
rect 1783 541 1967 575
rect 2025 677 2143 695
rect 2025 643 2109 677
rect 2025 609 2143 643
rect 2025 575 2109 609
rect 2025 559 2143 575
rect 1419 499 1967 541
rect 775 483 1158 495
rect 775 449 783 483
rect 817 479 1158 483
rect 817 449 972 479
rect 775 445 972 449
rect 1006 445 1040 479
rect 1074 445 1108 479
rect 1142 445 1158 479
rect 775 433 1158 445
rect 896 429 1158 433
rect 1192 429 1570 465
rect 595 391 862 399
rect 595 357 744 391
rect 778 357 812 391
rect 846 357 862 391
rect 595 349 862 357
rect 595 299 653 349
rect 896 315 962 429
rect 1192 395 1258 429
rect 1504 395 1570 429
rect 595 265 611 299
rect 645 265 653 299
rect 595 197 653 265
rect 595 163 611 197
rect 645 163 653 197
rect 595 147 653 163
rect 687 299 741 315
rect 687 265 697 299
rect 731 265 741 299
rect 687 193 741 265
rect 687 159 697 193
rect 731 159 741 193
rect 687 119 741 159
rect 775 299 962 315
rect 775 265 783 299
rect 817 265 962 299
rect 775 249 962 265
rect 1010 361 1052 395
rect 1086 361 1128 395
rect 1010 315 1128 361
rect 1010 281 1052 315
rect 1086 281 1128 315
rect 775 197 837 249
rect 775 163 783 197
rect 817 163 837 197
rect 775 147 837 163
rect 1010 233 1128 281
rect 1010 199 1052 233
rect 1086 199 1128 233
rect 1010 153 1128 199
rect 687 113 697 119
rect 619 107 697 113
rect 619 73 625 107
rect 659 85 697 107
rect 731 113 741 119
rect 1010 119 1052 153
rect 1086 119 1128 153
rect 1192 361 1208 395
rect 1242 361 1258 395
rect 1192 315 1258 361
rect 1192 281 1208 315
rect 1242 281 1258 315
rect 1192 233 1258 281
rect 1192 199 1208 233
rect 1242 199 1258 233
rect 1192 153 1258 199
rect 1192 119 1208 153
rect 1242 119 1258 153
rect 1322 361 1364 395
rect 1398 361 1440 395
rect 1322 315 1440 361
rect 1322 281 1364 315
rect 1398 281 1440 315
rect 1322 233 1440 281
rect 1322 199 1364 233
rect 1398 199 1440 233
rect 1322 153 1440 199
rect 1322 119 1364 153
rect 1398 119 1440 153
rect 731 107 809 113
rect 731 85 769 107
rect 659 73 769 85
rect 803 73 809 107
rect 619 67 809 73
rect 1010 85 1016 119
rect 1050 85 1088 119
rect 1122 85 1128 119
rect 1322 85 1328 119
rect 1362 85 1400 119
rect 1434 85 1440 119
rect 1010 51 1440 85
rect 1504 361 1520 395
rect 1554 361 1570 395
rect 1504 315 1570 361
rect 1504 281 1520 315
rect 1554 281 1570 315
rect 1504 233 1570 281
rect 1504 199 1520 233
rect 1554 199 1570 233
rect 1504 153 1570 199
rect 1504 119 1520 153
rect 1554 119 1570 153
rect 1634 395 1752 499
rect 1634 361 1676 395
rect 1710 361 1752 395
rect 1634 315 1752 361
rect 1634 281 1676 315
rect 1710 281 1752 315
rect 1634 233 1752 281
rect 1634 199 1676 233
rect 1710 199 1752 233
rect 1634 153 1752 199
rect 1634 119 1676 153
rect 1710 119 1752 153
rect 1816 395 1882 411
rect 1816 361 1832 395
rect 1866 361 1882 395
rect 1816 315 1882 361
rect 1816 281 1832 315
rect 1866 281 1882 315
rect 1816 233 1882 281
rect 1816 199 1832 233
rect 1866 199 1882 233
rect 1816 153 1882 199
rect 1816 119 1832 153
rect 1866 119 1882 153
rect 1504 85 1570 119
rect 1816 85 1882 119
rect 1504 51 1882 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 635 1509 669 1543
rect 707 1509 741 1543
rect 947 1509 981 1543
rect 1019 1509 1053 1543
rect 1944 1509 1978 1543
rect 2016 1509 2050 1543
rect 31 797 65 831
rect 1484 899 1518 933
rect 1556 899 1590 933
rect 1944 899 1978 933
rect 2016 899 2050 933
rect 697 610 731 644
rect 769 621 803 655
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 1597 695 1631 729
rect 1669 695 1703 729
rect 2031 695 2065 729
rect 2103 695 2137 729
rect 625 73 659 107
rect 697 85 731 119
rect 769 73 803 107
rect 1016 85 1050 119
rect 1088 85 1122 119
rect 1328 85 1362 119
rect 1400 85 1434 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 1645 2208 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2208 1645
rect 0 1605 2208 1611
rect 0 1543 2208 1577
rect 0 1509 635 1543
rect 669 1509 707 1543
rect 741 1509 947 1543
rect 981 1509 1019 1543
rect 1053 1509 1944 1543
rect 1978 1509 2016 1543
rect 2050 1509 2208 1543
rect 0 1503 2208 1509
rect 0 933 2208 939
rect 0 899 1484 933
rect 1518 899 1556 933
rect 1590 899 1944 933
rect 1978 899 2016 933
rect 2050 899 2208 933
rect 0 865 2208 899
rect 0 831 2208 837
rect 0 797 31 831
rect 65 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2208 831
rect 0 791 2208 797
rect 0 729 2208 763
rect 0 695 1597 729
rect 1631 695 1669 729
rect 1703 695 2031 729
rect 2065 695 2103 729
rect 2137 695 2208 729
rect 0 689 2208 695
rect 14 655 2194 661
rect 14 644 769 655
rect 14 610 697 644
rect 731 621 769 644
rect 803 621 2194 655
rect 731 610 2194 621
rect 14 604 2194 610
rect 0 119 2208 125
rect 0 107 697 119
rect 0 73 625 107
rect 659 85 697 107
rect 731 107 1016 119
rect 731 85 769 107
rect 659 73 769 85
rect 803 85 1016 107
rect 1050 85 1088 119
rect 1122 85 1328 119
rect 1362 85 1400 119
rect 1434 85 2208 119
rect 803 73 2208 85
rect 0 51 2208 73
rect 0 17 2208 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -23 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 lsbuflv2hv_1
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2143 1204 2177 1238 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2143 1130 2177 1164 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2143 1056 2177 1090 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2143 1278 2177 1312 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2143 1352 2177 1386 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel metal1 s 0 689 2208 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 865 2208 939 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 14 604 2194 661 0 FreeSans 340 0 0 0 LVPWR
port 2 nsew power bidirectional
flabel metal1 s 0 1605 2208 1628 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 0 2208 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 1503 2208 1577 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 51 2208 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 791 2208 837 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
rlabel viali s 769 621 803 655 1 LVPWR
port 2 nsew power bidirectional
rlabel viali s 697 610 731 644 1 LVPWR
port 2 nsew power bidirectional
rlabel metal1 s 14 604 2194 661 1 LVPWR
port 2 nsew power bidirectional
rlabel locali s 941 1233 1059 1543 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 629 1543 1059 1577 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 629 1233 747 1543 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1322 85 1440 395 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1010 85 1128 395 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1010 51 1440 85 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1938 1367 2056 1549 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 2016 1509 2050 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1944 1509 1978 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1400 85 1434 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1328 85 1362 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1088 85 1122 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1019 1509 1053 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1016 85 1050 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 947 1509 981 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 769 73 803 107 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 707 1509 741 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 697 85 731 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 635 1509 669 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 625 73 659 107 1 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 51 2208 125 1 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 1503 2208 1577 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 0 1611 2208 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 2143 1611 2177 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 2143 -17 2177 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 2047 1611 2081 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 2047 -17 2081 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1951 1611 1985 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1951 -17 1985 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1855 1611 1889 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1855 -17 1889 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1759 1611 1793 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1759 -17 1793 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1663 1611 1697 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1663 -17 1697 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1567 1611 1601 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1471 1611 1505 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1375 1611 1409 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1279 1611 1313 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1183 1611 1217 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1087 1611 1121 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 991 1611 1025 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 895 1611 929 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 895 -17 929 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 799 1611 833 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 799 -17 833 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 703 1611 737 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 703 -17 737 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 607 1611 641 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 607 -17 641 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 511 1611 545 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 511 -17 545 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 415 1611 449 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 415 -17 449 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 319 1611 353 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 319 -17 353 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 223 1611 257 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 223 -17 257 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 127 1611 161 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 127 -17 161 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 31 1611 65 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 31 -17 65 17 1 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 2208 23 1 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 1605 2208 1651 1 VNB
port 4 nsew ground bidirectional
rlabel locali s 1647 797 2208 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 2143 797 2177 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 2047 797 2081 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 1951 797 1985 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 1855 797 1889 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 1759 797 1793 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 1663 797 1697 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 31 797 65 831 1 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 791 2208 837 1 VPB
port 5 nsew power bidirectional
rlabel locali s 1478 881 1596 1189 1 VPWR
port 6 nsew power bidirectional
rlabel locali s 1591 575 1709 741 1 VPWR
port 6 nsew power bidirectional
rlabel locali s 1938 881 2056 1189 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 2103 695 2137 729 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 2031 695 2065 729 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 2016 899 2050 933 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1944 899 1978 933 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1669 695 1703 729 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1597 695 1631 729 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1556 899 1590 933 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1484 899 1518 933 1 VPWR
port 6 nsew power bidirectional
rlabel metal1 s 0 689 2208 763 1 VPWR
port 6 nsew power bidirectional
rlabel metal1 s 0 865 2208 939 1 VPWR
port 6 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 2208 1628
string GDS_END 272530
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 249164
string LEFclass CORE
string LEFsite unithvdbl
string LEFsymmetry X Y
<< end >>
