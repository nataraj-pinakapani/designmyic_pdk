magic
tech minimum
magscale 1 2
timestamp 1644097196
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 1 7 25 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 51 7 75 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 7 24 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 51 7 75 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 75 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 75 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 75 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 75 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 8 75 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 8 75 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 7 75 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 7 75 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 8 74 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 8 74 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 7 74 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 7 74 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 11 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 10 74 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 9 74 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 8 74 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 8 74 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 7 74 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 74 7 74 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 8 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 8 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 7 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 7 73 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 8 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 8 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 7 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 73 7 73 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 73 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 73 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 73 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 8 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 8 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 7 73 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 7 73 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 8 72 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 8 72 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 7 72 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 7 72 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 11 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 10 72 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 9 72 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 8 72 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 8 72 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 7 72 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 72 7 72 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 8 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 8 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 7 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 7 71 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 8 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 8 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 7 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 71 7 71 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 71 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 71 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 71 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 8 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 8 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 7 71 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 7 71 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 8 70 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 8 70 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 7 70 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 7 70 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 11 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 10 70 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 9 70 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 8 70 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 8 70 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 7 70 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 70 7 70 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 8 69 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 8 69 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 7 69 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 7 69 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 11 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 10 69 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 9 69 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 8 69 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 8 69 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 7 69 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 69 7 69 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 8 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 8 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 7 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 7 68 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 8 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 8 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 7 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 68 7 68 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 68 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 68 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 68 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 8 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 8 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 7 68 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 7 68 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 8 67 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 8 67 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 7 67 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 7 67 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 11 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 10 67 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 9 67 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 8 67 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 8 67 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 7 67 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 67 7 67 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 8 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 8 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 7 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 7 66 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 8 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 8 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 7 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 66 7 66 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 66 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 66 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 66 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 8 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 8 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 7 66 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 7 66 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 8 65 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 8 65 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 7 65 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 7 65 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 11 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 10 65 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 9 65 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 8 65 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 8 65 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 7 65 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 65 7 65 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 8 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 8 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 7 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 7 64 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 8 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 8 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 7 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 64 7 64 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 64 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 64 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 64 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 8 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 8 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 7 64 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 7 64 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 8 63 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 8 63 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 7 63 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 7 63 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 11 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 10 63 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 9 63 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 8 63 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 8 63 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 7 63 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 63 7 63 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 8 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 8 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 7 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 7 62 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 8 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 8 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 7 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 62 7 62 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 62 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 62 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 62 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 8 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 8 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 7 62 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 7 62 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 8 61 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 8 61 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 7 61 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 7 61 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 11 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 10 61 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 9 61 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 8 61 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 8 61 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 7 61 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 61 7 61 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 8 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 8 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 7 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 7 60 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 8 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 8 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 7 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 60 7 60 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 60 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 60 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 60 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 8 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 8 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 7 60 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 7 60 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 8 59 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 8 59 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 7 59 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 7 59 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 11 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 10 59 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 9 59 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 8 59 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 8 59 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 7 59 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 59 7 59 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 8 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 8 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 7 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 7 58 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 8 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 8 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 7 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 58 7 58 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 58 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 58 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 58 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 8 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 8 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 7 58 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 7 58 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 8 57 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 8 57 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 7 57 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 7 57 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 11 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 10 57 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 9 57 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 8 57 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 8 57 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 7 57 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 57 7 57 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 8 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 8 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 7 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 7 56 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 8 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 8 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 7 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 56 7 56 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 56 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 56 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 56 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 8 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 8 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 7 56 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 7 56 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 8 55 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 8 55 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 7 55 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 7 55 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 11 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 10 55 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 9 55 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 8 55 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 8 55 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 7 55 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 55 7 55 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 8 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 8 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 7 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 7 54 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 8 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 8 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 7 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 54 7 54 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 54 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 54 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 54 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 8 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 8 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 7 54 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 7 54 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 53 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 9 53 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 8 53 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 8 53 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 7 53 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 53 7 53 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 53 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 53 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 53 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 53 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 8 53 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 8 53 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 7 53 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 7 53 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 8 52 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 8 52 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 7 52 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 7 52 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 11 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 10 52 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 9 52 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 8 52 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 8 52 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 7 52 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 52 7 52 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 51 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 51 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 8 51 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 8 51 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 7 51 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 7 51 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 11 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 10 51 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 51 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 9 51 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 8 51 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 8 51 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 7 51 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 51 7 51 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 8 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 8 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 7 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 7 24 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 8 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 8 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 7 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 24 7 24 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 24 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 24 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 24 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 8 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 8 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 7 24 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 7 24 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 8 23 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 8 23 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 7 23 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 7 23 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 11 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 10 23 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 9 23 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 8 23 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 8 23 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 7 23 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 23 7 23 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 8 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 8 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 7 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 7 22 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 8 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 8 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 7 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 22 7 22 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 22 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 22 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 22 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 8 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 8 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 7 22 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 7 22 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 8 21 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 8 21 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 7 21 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 7 21 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 11 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 10 21 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 9 21 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 8 21 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 8 21 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 7 21 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 21 7 21 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 8 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 8 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 7 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 7 20 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 8 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 8 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 7 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 20 7 20 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 20 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 20 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 20 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 8 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 8 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 7 20 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 7 20 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 8 19 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 8 19 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 7 19 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 7 19 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 11 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 10 19 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 9 19 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 8 19 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 8 19 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 7 19 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 19 7 19 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 8 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 8 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 7 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 7 18 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 8 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 8 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 7 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 18 7 18 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 18 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 18 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 18 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 8 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 8 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 7 18 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 7 18 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 8 17 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 8 17 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 7 17 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 7 17 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 11 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 10 17 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 9 17 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 8 17 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 8 17 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 7 17 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 17 7 17 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 8 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 8 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 7 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 7 16 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 8 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 8 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 7 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 16 7 16 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 16 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 16 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 16 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 8 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 8 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 7 16 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 7 16 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 15 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 9 15 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 8 15 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 8 15 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 7 15 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 15 7 15 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 15 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 15 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 15 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 15 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 8 15 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 8 15 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 7 15 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 7 15 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 8 14 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 8 14 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 7 14 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 7 14 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 11 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 10 14 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 9 14 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 8 14 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 8 14 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 7 14 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 14 7 14 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 8 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 8 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 7 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 7 13 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 8 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 8 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 7 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 13 7 13 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 13 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 13 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 13 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 8 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 8 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 7 13 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 7 13 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 8 12 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 8 12 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 7 12 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 7 12 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 11 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 10 12 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 9 12 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 8 12 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 8 12 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 7 12 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 12 7 12 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 8 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 8 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 7 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 7 11 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 8 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 8 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 7 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 11 7 11 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 11 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 11 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 11 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 8 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 8 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 7 11 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 7 11 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 8 10 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 8 10 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 7 10 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 7 10 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 11 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 10 10 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 9 10 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 8 10 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 8 10 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 7 10 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 10 7 10 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 8 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 8 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 7 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 7 9 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 8 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 8 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 7 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 9 7 9 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 9 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 9 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 9 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 8 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 8 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 7 9 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 7 9 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 8 8 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 8 8 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 7 8 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 7 8 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 11 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 10 8 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 9 8 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 8 8 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 8 8 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 7 8 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 8 7 8 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 8 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 8 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 7 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 7 7 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 8 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 8 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 7 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 7 7 7 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 7 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 7 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 7 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 8 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 8 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 7 7 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 7 7 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 8 6 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 8 6 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 7 6 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 7 6 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 11 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 10 6 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 9 6 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 8 6 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 8 6 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 7 6 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 6 7 6 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 8 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 8 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 7 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 7 5 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 8 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 8 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 7 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 5 7 5 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 5 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 5 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 5 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 8 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 8 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 7 5 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 7 5 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 8 4 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 8 4 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 7 4 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 7 4 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 11 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 10 4 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 9 4 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 8 4 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 8 4 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 7 4 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 4 7 4 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 8 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 8 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 7 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 7 3 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 8 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 8 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 7 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 3 7 3 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 3 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 3 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 3 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 8 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 8 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 7 3 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 7 3 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 8 2 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 8 2 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 7 2 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 7 2 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 11 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 10 2 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 9 2 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 8 2 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 8 2 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 7 2 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 2 7 2 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 8 1 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 8 1 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 7 1 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 7 1 7 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 11 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 11 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 10 1 10 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 9 1 9 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 8 1 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 8 1 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 7 1 8 6 VCCD
port 3 nsew power bidirectional
rlabel nfet_brown s 1 7 1 7 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 46 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 54 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 198
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
