magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< locali >>
rect 0 1420 54 1476
rect 1662 1456 1716 1504
rect 88 1445 1716 1456
rect 88 1422 1672 1445
rect 0 1386 10 1420
rect 44 1386 54 1420
rect 1662 1411 1672 1422
rect 1706 1411 1716 1445
rect 0 1352 1628 1386
rect 1662 1373 1716 1411
rect 0 1348 54 1352
rect 0 1314 10 1348
rect 44 1314 54 1348
rect 1662 1339 1672 1373
rect 1706 1339 1716 1373
rect 1662 1316 1716 1339
rect 0 1276 54 1314
rect 88 1301 1716 1316
rect 88 1282 1672 1301
rect 0 1242 10 1276
rect 44 1246 54 1276
rect 1662 1267 1672 1282
rect 1706 1267 1716 1301
rect 44 1242 1628 1246
rect 0 1212 1628 1242
rect 1662 1229 1716 1267
rect 0 1204 54 1212
rect 0 1170 10 1204
rect 44 1170 54 1204
rect 1662 1195 1672 1229
rect 1706 1195 1716 1229
rect 1662 1176 1716 1195
rect 0 1132 54 1170
rect 88 1157 1716 1176
rect 88 1142 1672 1157
rect 0 1098 10 1132
rect 44 1106 54 1132
rect 1662 1123 1672 1142
rect 1706 1123 1716 1157
rect 44 1098 1628 1106
rect 0 1072 1628 1098
rect 1662 1085 1716 1123
rect 0 1060 54 1072
rect 0 1026 10 1060
rect 44 1026 54 1060
rect 1662 1051 1672 1085
rect 1706 1051 1716 1085
rect 1662 1036 1716 1051
rect 0 988 54 1026
rect 88 1013 1716 1036
rect 88 1002 1672 1013
rect 0 954 10 988
rect 44 966 54 988
rect 1662 979 1672 1002
rect 1706 979 1716 1013
rect 44 954 1628 966
rect 0 932 1628 954
rect 1662 941 1716 979
rect 0 916 54 932
rect 0 882 10 916
rect 44 882 54 916
rect 1662 907 1672 941
rect 1706 907 1716 941
rect 1662 896 1716 907
rect 0 844 54 882
rect 88 869 1716 896
rect 88 862 1672 869
rect 0 810 10 844
rect 44 826 54 844
rect 1662 835 1672 862
rect 1706 835 1716 869
rect 44 810 1628 826
rect 0 792 1628 810
rect 1662 797 1716 835
rect 0 772 54 792
rect 0 738 10 772
rect 44 738 54 772
rect 1662 763 1672 797
rect 1706 763 1716 797
rect 1662 756 1716 763
rect 0 700 54 738
rect 88 725 1716 756
rect 88 722 1672 725
rect 0 666 10 700
rect 44 686 54 700
rect 1662 691 1672 722
rect 1706 691 1716 725
rect 44 666 1628 686
rect 0 652 1628 666
rect 1662 653 1716 691
rect 0 628 54 652
rect 0 594 10 628
rect 44 594 54 628
rect 1662 619 1672 653
rect 1706 619 1716 653
rect 1662 616 1716 619
rect 0 556 54 594
rect 88 582 1716 616
rect 0 522 10 556
rect 44 546 54 556
rect 1662 581 1716 582
rect 1662 547 1672 581
rect 1706 547 1716 581
rect 44 522 1628 546
rect 0 512 1628 522
rect 0 484 54 512
rect 0 450 10 484
rect 44 450 54 484
rect 1662 509 1716 547
rect 1662 476 1672 509
rect 0 412 54 450
rect 88 475 1672 476
rect 1706 475 1716 509
rect 88 442 1716 475
rect 0 378 10 412
rect 44 406 54 412
rect 1662 437 1716 442
rect 44 378 1628 406
rect 0 372 1628 378
rect 1662 403 1672 437
rect 1706 403 1716 437
rect 0 340 54 372
rect 0 306 10 340
rect 44 306 54 340
rect 1662 365 1716 403
rect 1662 336 1672 365
rect 0 268 54 306
rect 88 331 1672 336
rect 1706 331 1716 365
rect 88 302 1716 331
rect 0 234 10 268
rect 44 266 54 268
rect 1662 293 1716 302
rect 44 234 1628 266
rect 0 232 1628 234
rect 1662 259 1672 293
rect 1706 259 1716 293
rect 0 196 54 232
rect 1662 221 1716 259
rect 1662 196 1672 221
rect 0 162 10 196
rect 44 162 54 196
rect 88 187 1672 196
rect 1706 187 1716 221
rect 88 162 1716 187
rect 0 126 54 162
rect 1662 149 1716 162
rect 0 124 1628 126
rect 0 90 10 124
rect 44 92 1628 124
rect 1662 115 1672 149
rect 1706 115 1716 149
rect 1662 92 1716 115
rect 44 90 54 92
rect 0 64 54 90
<< viali >>
rect 10 1386 44 1420
rect 1672 1411 1706 1445
rect 10 1314 44 1348
rect 1672 1339 1706 1373
rect 10 1242 44 1276
rect 1672 1267 1706 1301
rect 10 1170 44 1204
rect 1672 1195 1706 1229
rect 10 1098 44 1132
rect 1672 1123 1706 1157
rect 10 1026 44 1060
rect 1672 1051 1706 1085
rect 10 954 44 988
rect 1672 979 1706 1013
rect 10 882 44 916
rect 1672 907 1706 941
rect 10 810 44 844
rect 1672 835 1706 869
rect 10 738 44 772
rect 1672 763 1706 797
rect 10 666 44 700
rect 1672 691 1706 725
rect 10 594 44 628
rect 1672 619 1706 653
rect 10 522 44 556
rect 1672 547 1706 581
rect 10 450 44 484
rect 1672 475 1706 509
rect 10 378 44 412
rect 1672 403 1706 437
rect 10 306 44 340
rect 1672 331 1706 365
rect 10 234 44 268
rect 1672 259 1706 293
rect 10 162 44 196
rect 1672 187 1706 221
rect 10 90 44 124
rect 1672 115 1706 149
<< metal1 >>
rect 0 1562 1716 1568
rect 0 1510 76 1562
rect 128 1510 140 1562
rect 192 1510 204 1562
rect 256 1510 268 1562
rect 320 1510 332 1562
rect 384 1510 396 1562
rect 448 1510 460 1562
rect 512 1510 524 1562
rect 576 1510 588 1562
rect 640 1510 652 1562
rect 704 1510 716 1562
rect 768 1510 780 1562
rect 832 1510 844 1562
rect 896 1510 908 1562
rect 960 1510 972 1562
rect 1024 1510 1036 1562
rect 1088 1510 1100 1562
rect 1152 1510 1164 1562
rect 1216 1510 1228 1562
rect 1280 1510 1292 1562
rect 1344 1510 1356 1562
rect 1408 1510 1420 1562
rect 1472 1510 1484 1562
rect 1536 1510 1548 1562
rect 1600 1510 1612 1562
rect 1664 1510 1716 1562
rect 0 1504 1716 1510
rect 0 1449 54 1476
rect 0 1397 1 1449
rect 53 1397 54 1449
rect 0 1386 10 1397
rect 44 1386 54 1397
rect 0 1385 54 1386
rect 0 1333 1 1385
rect 53 1333 54 1385
rect 0 1321 10 1333
rect 44 1321 54 1333
rect 0 1269 1 1321
rect 53 1269 54 1321
rect 0 1257 10 1269
rect 44 1257 54 1269
rect 0 1205 1 1257
rect 53 1205 54 1257
rect 0 1204 54 1205
rect 0 1193 10 1204
rect 44 1193 54 1204
rect 0 1141 1 1193
rect 53 1141 54 1193
rect 0 1132 54 1141
rect 0 1129 10 1132
rect 44 1129 54 1132
rect 0 1077 1 1129
rect 53 1077 54 1129
rect 0 1065 54 1077
rect 0 1013 1 1065
rect 53 1013 54 1065
rect 0 1001 54 1013
rect 0 949 1 1001
rect 53 949 54 1001
rect 0 937 54 949
rect 0 885 1 937
rect 53 885 54 937
rect 0 882 10 885
rect 44 882 54 885
rect 0 873 54 882
rect 0 821 1 873
rect 53 821 54 873
rect 0 810 10 821
rect 44 810 54 821
rect 0 809 54 810
rect 0 757 1 809
rect 53 757 54 809
rect 0 745 10 757
rect 44 745 54 757
rect 0 693 1 745
rect 53 693 54 745
rect 0 681 10 693
rect 44 681 54 693
rect 0 629 1 681
rect 53 629 54 681
rect 0 628 54 629
rect 0 617 10 628
rect 44 617 54 628
rect 0 565 1 617
rect 53 565 54 617
rect 0 556 54 565
rect 0 553 10 556
rect 44 553 54 556
rect 0 501 1 553
rect 53 501 54 553
rect 0 489 54 501
rect 0 437 1 489
rect 53 437 54 489
rect 0 425 54 437
rect 0 373 1 425
rect 53 373 54 425
rect 0 361 54 373
rect 0 309 1 361
rect 53 309 54 361
rect 0 306 10 309
rect 44 306 54 309
rect 0 297 54 306
rect 0 245 1 297
rect 53 245 54 297
rect 0 234 10 245
rect 44 234 54 245
rect 0 233 54 234
rect 0 181 1 233
rect 53 181 54 233
rect 0 169 10 181
rect 44 169 54 181
rect 0 117 1 169
rect 53 117 54 169
rect 0 105 10 117
rect 44 105 54 117
rect 0 53 1 105
rect 53 64 54 105
rect 88 64 116 1476
rect 144 92 172 1504
rect 200 64 228 1476
rect 256 92 284 1504
rect 312 64 340 1476
rect 368 92 396 1504
rect 424 64 452 1476
rect 480 92 508 1504
rect 536 64 564 1476
rect 592 92 620 1504
rect 648 64 676 1476
rect 704 92 732 1504
rect 760 64 788 1476
rect 816 92 844 1504
rect 872 64 900 1476
rect 928 92 956 1504
rect 984 64 1012 1476
rect 1040 92 1068 1504
rect 1096 64 1124 1476
rect 1152 92 1180 1504
rect 1208 64 1236 1476
rect 1264 92 1292 1504
rect 1320 64 1348 1476
rect 1376 92 1404 1504
rect 1432 64 1460 1476
rect 1488 92 1516 1504
rect 1544 64 1572 1476
rect 1600 92 1628 1504
rect 1662 1494 1716 1504
rect 1662 1442 1663 1494
rect 1715 1442 1716 1494
rect 1662 1430 1672 1442
rect 1706 1430 1716 1442
rect 1662 1378 1663 1430
rect 1715 1378 1716 1430
rect 1662 1373 1716 1378
rect 1662 1366 1672 1373
rect 1706 1366 1716 1373
rect 1662 1314 1663 1366
rect 1715 1314 1716 1366
rect 1662 1302 1716 1314
rect 1662 1250 1663 1302
rect 1715 1250 1716 1302
rect 1662 1238 1716 1250
rect 1662 1186 1663 1238
rect 1715 1186 1716 1238
rect 1662 1174 1716 1186
rect 1662 1122 1663 1174
rect 1715 1122 1716 1174
rect 1662 1110 1716 1122
rect 1662 1058 1663 1110
rect 1715 1058 1716 1110
rect 1662 1051 1672 1058
rect 1706 1051 1716 1058
rect 1662 1046 1716 1051
rect 1662 994 1663 1046
rect 1715 994 1716 1046
rect 1662 982 1672 994
rect 1706 982 1716 994
rect 1662 930 1663 982
rect 1715 930 1716 982
rect 1662 918 1672 930
rect 1706 918 1716 930
rect 1662 866 1663 918
rect 1715 866 1716 918
rect 1662 854 1672 866
rect 1706 854 1716 866
rect 1662 802 1663 854
rect 1715 802 1716 854
rect 1662 797 1716 802
rect 1662 790 1672 797
rect 1706 790 1716 797
rect 1662 738 1663 790
rect 1715 738 1716 790
rect 1662 726 1716 738
rect 1662 674 1663 726
rect 1715 674 1716 726
rect 1662 662 1716 674
rect 1662 610 1663 662
rect 1715 610 1716 662
rect 1662 598 1716 610
rect 1662 546 1663 598
rect 1715 546 1716 598
rect 1662 534 1716 546
rect 1662 482 1663 534
rect 1715 482 1716 534
rect 1662 475 1672 482
rect 1706 475 1716 482
rect 1662 470 1716 475
rect 1662 418 1663 470
rect 1715 418 1716 470
rect 1662 406 1672 418
rect 1706 406 1716 418
rect 1662 354 1663 406
rect 1715 354 1716 406
rect 1662 342 1672 354
rect 1706 342 1716 354
rect 1662 290 1663 342
rect 1715 290 1716 342
rect 1662 278 1672 290
rect 1706 278 1716 290
rect 1662 226 1663 278
rect 1715 226 1716 278
rect 1662 221 1716 226
rect 1662 214 1672 221
rect 1706 214 1716 221
rect 1662 162 1663 214
rect 1715 162 1716 214
rect 1662 150 1716 162
rect 1662 98 1663 150
rect 1715 98 1716 150
rect 1662 92 1716 98
rect 53 58 1716 64
rect 53 53 76 58
rect 0 6 76 53
rect 128 6 140 58
rect 192 6 204 58
rect 256 6 268 58
rect 320 6 332 58
rect 384 6 396 58
rect 448 6 460 58
rect 512 6 524 58
rect 576 6 588 58
rect 640 6 652 58
rect 704 6 716 58
rect 768 6 780 58
rect 832 6 844 58
rect 896 6 908 58
rect 960 6 972 58
rect 1024 6 1036 58
rect 1088 6 1100 58
rect 1152 6 1164 58
rect 1216 6 1228 58
rect 1280 6 1292 58
rect 1344 6 1356 58
rect 1408 6 1420 58
rect 1472 6 1484 58
rect 1536 6 1548 58
rect 1600 6 1612 58
rect 1664 6 1716 58
rect 0 0 1716 6
<< via1 >>
rect 76 1510 128 1562
rect 140 1510 192 1562
rect 204 1510 256 1562
rect 268 1510 320 1562
rect 332 1510 384 1562
rect 396 1510 448 1562
rect 460 1510 512 1562
rect 524 1510 576 1562
rect 588 1510 640 1562
rect 652 1510 704 1562
rect 716 1510 768 1562
rect 780 1510 832 1562
rect 844 1510 896 1562
rect 908 1510 960 1562
rect 972 1510 1024 1562
rect 1036 1510 1088 1562
rect 1100 1510 1152 1562
rect 1164 1510 1216 1562
rect 1228 1510 1280 1562
rect 1292 1510 1344 1562
rect 1356 1510 1408 1562
rect 1420 1510 1472 1562
rect 1484 1510 1536 1562
rect 1548 1510 1600 1562
rect 1612 1510 1664 1562
rect 1 1420 53 1449
rect 1 1397 10 1420
rect 10 1397 44 1420
rect 44 1397 53 1420
rect 1 1348 53 1385
rect 1 1333 10 1348
rect 10 1333 44 1348
rect 44 1333 53 1348
rect 1 1314 10 1321
rect 10 1314 44 1321
rect 44 1314 53 1321
rect 1 1276 53 1314
rect 1 1269 10 1276
rect 10 1269 44 1276
rect 44 1269 53 1276
rect 1 1242 10 1257
rect 10 1242 44 1257
rect 44 1242 53 1257
rect 1 1205 53 1242
rect 1 1170 10 1193
rect 10 1170 44 1193
rect 44 1170 53 1193
rect 1 1141 53 1170
rect 1 1098 10 1129
rect 10 1098 44 1129
rect 44 1098 53 1129
rect 1 1077 53 1098
rect 1 1060 53 1065
rect 1 1026 10 1060
rect 10 1026 44 1060
rect 44 1026 53 1060
rect 1 1013 53 1026
rect 1 988 53 1001
rect 1 954 10 988
rect 10 954 44 988
rect 44 954 53 988
rect 1 949 53 954
rect 1 916 53 937
rect 1 885 10 916
rect 10 885 44 916
rect 44 885 53 916
rect 1 844 53 873
rect 1 821 10 844
rect 10 821 44 844
rect 44 821 53 844
rect 1 772 53 809
rect 1 757 10 772
rect 10 757 44 772
rect 44 757 53 772
rect 1 738 10 745
rect 10 738 44 745
rect 44 738 53 745
rect 1 700 53 738
rect 1 693 10 700
rect 10 693 44 700
rect 44 693 53 700
rect 1 666 10 681
rect 10 666 44 681
rect 44 666 53 681
rect 1 629 53 666
rect 1 594 10 617
rect 10 594 44 617
rect 44 594 53 617
rect 1 565 53 594
rect 1 522 10 553
rect 10 522 44 553
rect 44 522 53 553
rect 1 501 53 522
rect 1 484 53 489
rect 1 450 10 484
rect 10 450 44 484
rect 44 450 53 484
rect 1 437 53 450
rect 1 412 53 425
rect 1 378 10 412
rect 10 378 44 412
rect 44 378 53 412
rect 1 373 53 378
rect 1 340 53 361
rect 1 309 10 340
rect 10 309 44 340
rect 44 309 53 340
rect 1 268 53 297
rect 1 245 10 268
rect 10 245 44 268
rect 44 245 53 268
rect 1 196 53 233
rect 1 181 10 196
rect 10 181 44 196
rect 44 181 53 196
rect 1 162 10 169
rect 10 162 44 169
rect 44 162 53 169
rect 1 124 53 162
rect 1 117 10 124
rect 10 117 44 124
rect 44 117 53 124
rect 1 90 10 105
rect 10 90 44 105
rect 44 90 53 105
rect 1 53 53 90
rect 1663 1445 1715 1494
rect 1663 1442 1672 1445
rect 1672 1442 1706 1445
rect 1706 1442 1715 1445
rect 1663 1411 1672 1430
rect 1672 1411 1706 1430
rect 1706 1411 1715 1430
rect 1663 1378 1715 1411
rect 1663 1339 1672 1366
rect 1672 1339 1706 1366
rect 1706 1339 1715 1366
rect 1663 1314 1715 1339
rect 1663 1301 1715 1302
rect 1663 1267 1672 1301
rect 1672 1267 1706 1301
rect 1706 1267 1715 1301
rect 1663 1250 1715 1267
rect 1663 1229 1715 1238
rect 1663 1195 1672 1229
rect 1672 1195 1706 1229
rect 1706 1195 1715 1229
rect 1663 1186 1715 1195
rect 1663 1157 1715 1174
rect 1663 1123 1672 1157
rect 1672 1123 1706 1157
rect 1706 1123 1715 1157
rect 1663 1122 1715 1123
rect 1663 1085 1715 1110
rect 1663 1058 1672 1085
rect 1672 1058 1706 1085
rect 1706 1058 1715 1085
rect 1663 1013 1715 1046
rect 1663 994 1672 1013
rect 1672 994 1706 1013
rect 1706 994 1715 1013
rect 1663 979 1672 982
rect 1672 979 1706 982
rect 1706 979 1715 982
rect 1663 941 1715 979
rect 1663 930 1672 941
rect 1672 930 1706 941
rect 1706 930 1715 941
rect 1663 907 1672 918
rect 1672 907 1706 918
rect 1706 907 1715 918
rect 1663 869 1715 907
rect 1663 866 1672 869
rect 1672 866 1706 869
rect 1706 866 1715 869
rect 1663 835 1672 854
rect 1672 835 1706 854
rect 1706 835 1715 854
rect 1663 802 1715 835
rect 1663 763 1672 790
rect 1672 763 1706 790
rect 1706 763 1715 790
rect 1663 738 1715 763
rect 1663 725 1715 726
rect 1663 691 1672 725
rect 1672 691 1706 725
rect 1706 691 1715 725
rect 1663 674 1715 691
rect 1663 653 1715 662
rect 1663 619 1672 653
rect 1672 619 1706 653
rect 1706 619 1715 653
rect 1663 610 1715 619
rect 1663 581 1715 598
rect 1663 547 1672 581
rect 1672 547 1706 581
rect 1706 547 1715 581
rect 1663 546 1715 547
rect 1663 509 1715 534
rect 1663 482 1672 509
rect 1672 482 1706 509
rect 1706 482 1715 509
rect 1663 437 1715 470
rect 1663 418 1672 437
rect 1672 418 1706 437
rect 1706 418 1715 437
rect 1663 403 1672 406
rect 1672 403 1706 406
rect 1706 403 1715 406
rect 1663 365 1715 403
rect 1663 354 1672 365
rect 1672 354 1706 365
rect 1706 354 1715 365
rect 1663 331 1672 342
rect 1672 331 1706 342
rect 1706 331 1715 342
rect 1663 293 1715 331
rect 1663 290 1672 293
rect 1672 290 1706 293
rect 1706 290 1715 293
rect 1663 259 1672 278
rect 1672 259 1706 278
rect 1706 259 1715 278
rect 1663 226 1715 259
rect 1663 187 1672 214
rect 1672 187 1706 214
rect 1706 187 1715 214
rect 1663 162 1715 187
rect 1663 149 1715 150
rect 1663 115 1672 149
rect 1672 115 1706 149
rect 1706 115 1715 149
rect 1663 98 1715 115
rect 76 6 128 58
rect 140 6 192 58
rect 204 6 256 58
rect 268 6 320 58
rect 332 6 384 58
rect 396 6 448 58
rect 460 6 512 58
rect 524 6 576 58
rect 588 6 640 58
rect 652 6 704 58
rect 716 6 768 58
rect 780 6 832 58
rect 844 6 896 58
rect 908 6 960 58
rect 972 6 1024 58
rect 1036 6 1088 58
rect 1100 6 1152 58
rect 1164 6 1216 58
rect 1228 6 1280 58
rect 1292 6 1344 58
rect 1356 6 1408 58
rect 1420 6 1472 58
rect 1484 6 1536 58
rect 1548 6 1600 58
rect 1612 6 1664 58
<< metal2 >>
rect 0 1562 1716 1568
rect 0 1510 76 1562
rect 128 1510 140 1562
rect 192 1510 204 1562
rect 256 1510 268 1562
rect 320 1510 332 1562
rect 384 1510 396 1562
rect 448 1510 460 1562
rect 512 1510 524 1562
rect 576 1510 588 1562
rect 640 1510 652 1562
rect 704 1510 716 1562
rect 768 1510 780 1562
rect 832 1510 844 1562
rect 896 1510 908 1562
rect 960 1510 972 1562
rect 1024 1510 1036 1562
rect 1088 1510 1100 1562
rect 1152 1510 1164 1562
rect 1216 1510 1228 1562
rect 1280 1510 1292 1562
rect 1344 1510 1356 1562
rect 1408 1510 1420 1562
rect 1472 1510 1484 1562
rect 1536 1510 1548 1562
rect 1600 1510 1612 1562
rect 1664 1510 1716 1562
rect 0 1504 1716 1510
rect 0 1449 54 1476
rect 0 1397 1 1449
rect 53 1397 54 1449
rect 0 1385 54 1397
rect 0 1333 1 1385
rect 53 1333 54 1385
rect 0 1321 54 1333
rect 0 1269 1 1321
rect 53 1269 54 1321
rect 0 1257 54 1269
rect 0 1205 1 1257
rect 53 1205 54 1257
rect 0 1193 54 1205
rect 0 1141 1 1193
rect 53 1141 54 1193
rect 0 1129 54 1141
rect 0 1077 1 1129
rect 53 1077 54 1129
rect 0 1065 54 1077
rect 0 1013 1 1065
rect 53 1013 54 1065
rect 0 1001 54 1013
rect 0 949 1 1001
rect 53 949 54 1001
rect 0 937 54 949
rect 0 885 1 937
rect 53 885 54 937
rect 0 873 54 885
rect 0 821 1 873
rect 53 821 54 873
rect 0 809 54 821
rect 0 757 1 809
rect 53 757 54 809
rect 0 745 54 757
rect 0 693 1 745
rect 53 693 54 745
rect 0 681 54 693
rect 0 629 1 681
rect 53 629 54 681
rect 0 617 54 629
rect 0 565 1 617
rect 53 565 54 617
rect 0 553 54 565
rect 0 501 1 553
rect 53 501 54 553
rect 0 489 54 501
rect 0 437 1 489
rect 53 437 54 489
rect 0 425 54 437
rect 0 373 1 425
rect 53 373 54 425
rect 0 361 54 373
rect 0 309 1 361
rect 53 309 54 361
rect 0 297 54 309
rect 0 245 1 297
rect 53 245 54 297
rect 0 233 54 245
rect 0 181 1 233
rect 53 181 54 233
rect 0 169 54 181
rect 0 117 1 169
rect 53 117 54 169
rect 0 105 54 117
rect 0 53 1 105
rect 53 64 54 105
rect 88 92 116 1504
rect 144 64 172 1476
rect 200 92 228 1504
rect 256 64 284 1476
rect 312 92 340 1504
rect 368 64 396 1476
rect 424 92 452 1504
rect 480 64 508 1476
rect 536 92 564 1504
rect 592 64 620 1476
rect 648 92 676 1504
rect 704 64 732 1476
rect 760 92 788 1504
rect 816 64 844 1476
rect 872 92 900 1504
rect 928 64 956 1476
rect 984 92 1012 1504
rect 1040 64 1068 1476
rect 1096 92 1124 1504
rect 1152 64 1180 1476
rect 1208 92 1236 1504
rect 1264 64 1292 1476
rect 1320 92 1348 1504
rect 1376 64 1404 1476
rect 1432 92 1460 1504
rect 1488 64 1516 1476
rect 1544 92 1572 1504
rect 1662 1494 1716 1504
rect 1600 64 1628 1476
rect 1662 1442 1663 1494
rect 1715 1442 1716 1494
rect 1662 1430 1716 1442
rect 1662 1378 1663 1430
rect 1715 1378 1716 1430
rect 1662 1366 1716 1378
rect 1662 1314 1663 1366
rect 1715 1314 1716 1366
rect 1662 1302 1716 1314
rect 1662 1250 1663 1302
rect 1715 1250 1716 1302
rect 1662 1238 1716 1250
rect 1662 1186 1663 1238
rect 1715 1186 1716 1238
rect 1662 1174 1716 1186
rect 1662 1122 1663 1174
rect 1715 1122 1716 1174
rect 1662 1110 1716 1122
rect 1662 1058 1663 1110
rect 1715 1058 1716 1110
rect 1662 1046 1716 1058
rect 1662 994 1663 1046
rect 1715 994 1716 1046
rect 1662 982 1716 994
rect 1662 930 1663 982
rect 1715 930 1716 982
rect 1662 918 1716 930
rect 1662 866 1663 918
rect 1715 866 1716 918
rect 1662 854 1716 866
rect 1662 802 1663 854
rect 1715 802 1716 854
rect 1662 790 1716 802
rect 1662 738 1663 790
rect 1715 738 1716 790
rect 1662 726 1716 738
rect 1662 674 1663 726
rect 1715 674 1716 726
rect 1662 662 1716 674
rect 1662 610 1663 662
rect 1715 610 1716 662
rect 1662 598 1716 610
rect 1662 546 1663 598
rect 1715 546 1716 598
rect 1662 534 1716 546
rect 1662 482 1663 534
rect 1715 482 1716 534
rect 1662 470 1716 482
rect 1662 418 1663 470
rect 1715 418 1716 470
rect 1662 406 1716 418
rect 1662 354 1663 406
rect 1715 354 1716 406
rect 1662 342 1716 354
rect 1662 290 1663 342
rect 1715 290 1716 342
rect 1662 278 1716 290
rect 1662 226 1663 278
rect 1715 226 1716 278
rect 1662 214 1716 226
rect 1662 162 1663 214
rect 1715 162 1716 214
rect 1662 150 1716 162
rect 1662 98 1663 150
rect 1715 98 1716 150
rect 1662 92 1716 98
rect 53 58 1716 64
rect 53 53 76 58
rect 0 6 76 53
rect 128 6 140 58
rect 192 6 204 58
rect 256 6 268 58
rect 320 6 332 58
rect 384 6 396 58
rect 448 6 460 58
rect 512 6 524 58
rect 576 6 588 58
rect 640 6 652 58
rect 704 6 716 58
rect 768 6 780 58
rect 832 6 844 58
rect 896 6 908 58
rect 960 6 972 58
rect 1024 6 1036 58
rect 1088 6 1100 58
rect 1152 6 1164 58
rect 1216 6 1228 58
rect 1280 6 1292 58
rect 1344 6 1356 58
rect 1408 6 1420 58
rect 1472 6 1484 58
rect 1536 6 1548 58
rect 1600 6 1612 58
rect 1664 6 1716 58
rect 0 0 1716 6
<< properties >>
string GDS_END 256840
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 241220
<< end >>
