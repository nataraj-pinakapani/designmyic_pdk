magic
tech sky130B
timestamp 1663361622
<< properties >>
string GDS_END 3190980
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 3190464
<< end >>
