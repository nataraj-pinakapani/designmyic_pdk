magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 11 0 11 11 6 C0
port 1 nsew
rlabel  s 10 6 10 11 6 C0
port 1 nsew
rlabel  s 10 0 10 5 6 C0
port 1 nsew
rlabel  s 9 6 9 11 6 C0
port 1 nsew
rlabel  s 9 0 9 5 6 C0
port 1 nsew
rlabel  s 7 6 8 11 6 C0
port 1 nsew
rlabel  s 7 0 8 5 6 C0
port 1 nsew
rlabel  s 6 6 7 11 6 C0
port 1 nsew
rlabel  s 6 0 7 5 6 C0
port 1 nsew
rlabel  s 5 6 5 11 6 C0
port 1 nsew
rlabel  s 5 0 5 5 6 C0
port 1 nsew
rlabel  s 4 6 4 11 6 C0
port 1 nsew
rlabel  s 4 0 4 5 6 C0
port 1 nsew
rlabel  s 2 6 3 11 6 C0
port 1 nsew
rlabel  s 2 0 3 5 6 C0
port 1 nsew
rlabel  s 1 6 2 11 6 C0
port 1 nsew
rlabel  s 1 0 2 5 6 C0
port 1 nsew
rlabel  s 0 11 11 12 6 C0
port 1 nsew
rlabel  s 0 0 0 11 4 C0
port 1 nsew
rlabel  s 0 0 11 0 8 C0
port 1 nsew
rlabel  s 10 6 11 11 6 C1
port 2 nsew
rlabel  s 10 1 11 6 6 C1
port 2 nsew
rlabel  s 9 6 10 11 6 C1
port 2 nsew
rlabel  s 9 1 10 6 6 C1
port 2 nsew
rlabel  s 8 6 8 11 6 C1
port 2 nsew
rlabel  s 8 1 8 6 6 C1
port 2 nsew
rlabel  s 7 6 7 11 6 C1
port 2 nsew
rlabel  s 7 1 7 6 6 C1
port 2 nsew
rlabel  s 6 6 6 11 6 C1
port 2 nsew
rlabel  s 6 1 6 6 6 C1
port 2 nsew
rlabel  s 4 6 5 11 6 C1
port 2 nsew
rlabel  s 4 1 5 6 6 C1
port 2 nsew
rlabel  s 3 6 3 11 6 C1
port 2 nsew
rlabel  s 3 1 3 6 6 C1
port 2 nsew
rlabel  s 2 6 2 11 6 C1
port 2 nsew
rlabel  s 2 1 2 6 6 C1
port 2 nsew
rlabel  s 1 6 1 11 6 C1
port 2 nsew
rlabel  s 1 6 11 6 6 C1
port 2 nsew
rlabel  s 1 1 1 6 6 C1
port 2 nsew
rlabel metal_blue s 6 6 6 7 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 11 12
string LEFview TRUE
<< end >>
