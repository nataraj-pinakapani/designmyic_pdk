magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 546 897
<< pwell >>
rect 50 43 458 287
rect -26 -43 506 43
<< locali >>
rect 25 310 203 387
rect 244 339 294 751
rect 244 305 359 339
rect 395 305 455 371
rect 316 269 359 305
rect 316 235 436 269
rect 370 103 436 235
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 18 735 208 751
rect 18 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 208 735
rect 18 435 208 701
rect 332 735 450 751
rect 332 701 338 735
rect 372 701 410 735
rect 444 701 450 735
rect 332 435 450 701
rect 18 113 280 269
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 240 113
rect 274 79 280 113
rect 18 73 280 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 24 701 58 735
rect 96 701 130 735
rect 168 701 202 735
rect 338 701 372 735
rect 410 701 444 735
rect 24 79 58 113
rect 96 79 130 113
rect 168 79 202 113
rect 240 79 274 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 831 480 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 0 791 480 797
rect 0 735 480 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 338 735
rect 372 701 410 735
rect 444 701 480 735
rect 0 689 480 701
rect 0 113 480 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 240 113
rect 274 79 480 113
rect 0 51 480 79
rect 0 17 480 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -23 480 -17
<< labels >>
rlabel locali s 395 305 455 371 6 A
port 1 nsew signal input
rlabel locali s 25 310 203 387 6 B
port 2 nsew signal input
rlabel metal1 s 0 51 480 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 480 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 506 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 50 43 458 287 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 480 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 546 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 480 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 370 103 436 235 6 Y
port 7 nsew signal output
rlabel locali s 316 235 436 269 6 Y
port 7 nsew signal output
rlabel locali s 316 269 359 305 6 Y
port 7 nsew signal output
rlabel locali s 244 305 359 339 6 Y
port 7 nsew signal output
rlabel locali s 244 339 294 751 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 480 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 211558
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 204800
<< end >>
