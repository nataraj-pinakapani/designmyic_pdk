magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 3 3 3 5 6 DRAIN
port 1 nsew
rlabel  s 1 3 2 5 6 DRAIN
port 1 nsew
rlabel  s 0 5 4 8 6 DRAIN
port 1 nsew
rlabel  s 1 5 3 6 6 GATE
port 2 nsew
rlabel  s 1 2 3 2 6 GATE
port 2 nsew
rlabel  s 3 3 4 5 6 SOURCE
port 3 nsew
rlabel  s 2 3 3 5 6 SOURCE
port 3 nsew
rlabel  s 1 3 1 5 6 SOURCE
port 3 nsew
rlabel  s 0 0 4 3 6 SOURCE
port 3 nsew
rlabel  s 0 3 0 5 4 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 4 8
string LEFview TRUE
<< end >>
