magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel 
 s 17 0 19 1 8 PAD_A_ESD_H
port 1 nsew signal bidirectional
rlabel � s 17 0 19 1 8 PAD_A_ESD_H
port 1 nsew signal bidirectional
rlabel 
 s 29 0 30 0 8 XRES_H_N
port 2 nsew signal output
rlabel � s 29 0 30 0 8 XRES_H_N
port 2 nsew signal output
rlabel 
 s 20 0 21 1 8 FILT_IN_H
port 3 nsew signal input
rlabel � s 20 0 21 1 8 FILT_IN_H
port 3 nsew signal input
rlabel 
 s 8 0 9 0 8 ENABLE_VDDIO
port 4 nsew signal input
rlabel � s 8 0 9 0 8 ENABLE_VDDIO
port 4 nsew signal input
rlabel 
 s 72 0 73 0 8 TIE_WEAK_HI_H
port 5 nsew signal bidirectional
rlabel � s 72 0 73 0 8 TIE_WEAK_HI_H
port 5 nsew signal bidirectional
rlabel 
 s 72 50 74 64 6 TIE_WEAK_HI_H
port 5 nsew signal bidirectional
rlabel � s 12 0 13 0 8 ENABLE_H
port 6 nsew signal input
rlabel  s 12 0 13 0 8 ENABLE_H
port 6 nsew signal input
rlabel � s 15 0 15 0 8 PULLUP_H
port 7 nsew signal bidirectional
rlabel  s 15 0 15 0 8 PULLUP_H
port 7 nsew signal bidirectional
rlabel � s 22 0 23 0 8 EN_VDDIO_SIG_H
port 8 nsew signal input
rlabel  s 22 0 23 0 8 EN_VDDIO_SIG_H
port 8 nsew signal input
rlabel � s 29 5 30 11 6 EN_VDDIO_SIG_H
port 8 nsew signal input
rlabel � s 28 0 28 0 8 TIE_LO_ESD
port 9 nsew signal output
rlabel  s 28 0 28 0 8 TIE_LO_ESD
port 9 nsew signal output
rlabel � s 31 0 31 0 8 TIE_HI_ESD
port 10 nsew signal output
rlabel  s 31 0 31 0 8 TIE_HI_ESD
port 10 nsew signal output
rlabel � s 33 0 33 0 8 DISABLE_PULLUP_H
port 11 nsew signal input
rlabel  s 33 0 33 0 8 DISABLE_PULLUP_H
port 11 nsew signal input
rlabel  s 25 0 25 10 6 INP_SEL_H
port 12 nsew signal input
rlabel  s 0 176 1 200 4 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 13 nsew ground bidirectional
rlabel  s 0 176 1 200 4 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 26 75 30 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 176 75 200 6 VSSIO
port 13 nsew ground bidirectional
rlabel  s 0 26 1 30 4 VSSIO
port 13 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 14 nsew ground bidirectional
rlabel  s 0 56 75 57 6 VSSA
port 14 nsew ground bidirectional
rlabel  s 0 48 75 48 6 VSSA
port 14 nsew ground bidirectional
rlabel  s 74 52 75 53 6 VSSA
port 14 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 14 nsew ground bidirectional
rlabel  s 0 52 1 53 4 VSSA
port 14 nsew ground bidirectional
rlabel  s 74 48 75 57 6 VSSA
port 14 nsew ground bidirectional
rlabel  s 74 37 75 40 6 VSSA
port 14 nsew ground bidirectional
rlabel  s 0 37 1 40 4 VSSA
port 14 nsew ground bidirectional
rlabel  s 0 48 1 57 4 VSSA
port 14 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 15 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 15 nsew ground bidirectional
rlabel  s 74 42 75 46 6 VSSD
port 15 nsew ground bidirectional
rlabel  s 0 42 1 46 4 VSSD
port 15 nsew ground bidirectional
rlabel  s 0 48 75 51 6 AMUXBUS_B
port 16 nsew signal bidirectional
rlabel  s 0 53 75 56 6 AMUXBUS_A
port 17 nsew signal bidirectional
rlabel  s 74 64 75 69 6 VDDIO_Q
port 18 nsew power bidirectional
rlabel  s 0 64 1 69 4 VDDIO_Q
port 18 nsew power bidirectional
rlabel  s 74 64 75 68 6 VDDIO_Q
port 18 nsew power bidirectional
rlabel  s 0 64 1 68 4 VDDIO_Q
port 18 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 19 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 19 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 19 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 19 nsew power bidirectional
rlabel  s 74 20 75 24 6 VDDIO
port 19 nsew power bidirectional
rlabel  s 74 70 75 95 6 VDDIO
port 19 nsew power bidirectional
rlabel  s 0 70 1 95 4 VDDIO
port 19 nsew power bidirectional
rlabel  s 0 20 1 24 4 VDDIO
port 19 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 20 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 20 nsew power bidirectional
rlabel  s 74 32 75 35 6 VSWITCH
port 20 nsew power bidirectional
rlabel  s 0 32 1 35 4 VSWITCH
port 20 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 21 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 21 nsew power bidirectional
rlabel  s 74 15 75 18 6 VDDA
port 21 nsew power bidirectional
rlabel  s 0 15 1 18 4 VDDA
port 21 nsew power bidirectional
rlabel  s 74 9 75 14 6 VCCD
port 22 nsew power bidirectional
rlabel  s 0 9 1 14 4 VCCD
port 22 nsew power bidirectional
rlabel  s 74 9 75 13 6 VCCD
port 22 nsew power bidirectional
rlabel  s 0 9 1 13 4 VCCD
port 22 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 23 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 23 nsew power bidirectional
rlabel  s 74 2 75 7 6 VCCHIB
port 23 nsew power bidirectional
rlabel  s 0 2 1 7 4 VCCHIB
port 23 nsew power bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 24 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 24 nsew ground bidirectional
rlabel  s 74 58 75 63 6 VSSIO_Q
port 24 nsew ground bidirectional
rlabel  s 0 58 1 63 4 VSSIO_Q
port 24 nsew ground bidirectional
rlabel  s 17 108 54 164 6 PAD
port 25 nsew signal bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 200
string LEFsymmetry R90
string LEFview TRUE
<< end >>
