magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 21 43 727 283
rect -26 -43 794 43
<< mvnmos >>
rect 104 107 204 257
rect 246 107 346 257
rect 402 107 502 257
rect 544 107 644 257
<< mvpmos >>
rect 90 443 190 743
rect 246 443 346 743
rect 402 443 502 743
rect 558 443 658 743
<< mvndiff >>
rect 47 249 104 257
rect 47 215 59 249
rect 93 215 104 249
rect 47 149 104 215
rect 47 115 59 149
rect 93 115 104 149
rect 47 107 104 115
rect 204 107 246 257
rect 346 249 402 257
rect 346 215 357 249
rect 391 215 402 249
rect 346 149 402 215
rect 346 115 357 149
rect 391 115 402 149
rect 346 107 402 115
rect 502 107 544 257
rect 644 249 701 257
rect 644 215 655 249
rect 689 215 701 249
rect 644 149 701 215
rect 644 115 655 149
rect 689 115 701 149
rect 644 107 701 115
<< mvpdiff >>
rect 33 735 90 743
rect 33 701 45 735
rect 79 701 90 735
rect 33 652 90 701
rect 33 618 45 652
rect 79 618 90 652
rect 33 568 90 618
rect 33 534 45 568
rect 79 534 90 568
rect 33 485 90 534
rect 33 451 45 485
rect 79 451 90 485
rect 33 443 90 451
rect 190 691 246 743
rect 190 657 201 691
rect 235 657 246 691
rect 190 623 246 657
rect 190 589 201 623
rect 235 589 246 623
rect 190 553 246 589
rect 190 519 201 553
rect 235 519 246 553
rect 190 485 246 519
rect 190 451 201 485
rect 235 451 246 485
rect 190 443 246 451
rect 346 735 402 743
rect 346 701 357 735
rect 391 701 402 735
rect 346 652 402 701
rect 346 618 357 652
rect 391 618 402 652
rect 346 568 402 618
rect 346 534 357 568
rect 391 534 402 568
rect 346 485 402 534
rect 346 451 357 485
rect 391 451 402 485
rect 346 443 402 451
rect 502 735 558 743
rect 502 701 513 735
rect 547 701 558 735
rect 502 654 558 701
rect 502 620 513 654
rect 547 620 558 654
rect 502 571 558 620
rect 502 537 513 571
rect 547 537 558 571
rect 502 490 558 537
rect 502 456 513 490
rect 547 456 558 490
rect 502 443 558 456
rect 658 735 715 743
rect 658 701 669 735
rect 703 701 715 735
rect 658 652 715 701
rect 658 618 669 652
rect 703 618 715 652
rect 658 568 715 618
rect 658 534 669 568
rect 703 534 715 568
rect 658 485 715 534
rect 658 451 669 485
rect 703 451 715 485
rect 658 443 715 451
<< mvndiffc >>
rect 59 215 93 249
rect 59 115 93 149
rect 357 215 391 249
rect 357 115 391 149
rect 655 215 689 249
rect 655 115 689 149
<< mvpdiffc >>
rect 45 701 79 735
rect 45 618 79 652
rect 45 534 79 568
rect 45 451 79 485
rect 201 657 235 691
rect 201 589 235 623
rect 201 519 235 553
rect 201 451 235 485
rect 357 701 391 735
rect 357 618 391 652
rect 357 534 391 568
rect 357 451 391 485
rect 513 701 547 735
rect 513 620 547 654
rect 513 537 547 571
rect 513 456 547 490
rect 669 701 703 735
rect 669 618 703 652
rect 669 534 703 568
rect 669 451 703 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
<< poly >>
rect 90 743 190 769
rect 246 743 346 769
rect 402 743 502 769
rect 558 743 658 769
rect 90 417 190 443
rect 90 351 204 417
rect 90 317 110 351
rect 144 317 204 351
rect 90 283 204 317
rect 104 257 204 283
rect 246 383 346 443
rect 246 342 360 383
rect 246 308 309 342
rect 343 308 360 342
rect 246 283 360 308
rect 402 343 502 443
rect 558 417 658 443
rect 402 309 425 343
rect 459 309 502 343
rect 246 257 346 283
rect 402 257 502 309
rect 544 343 658 417
rect 544 309 604 343
rect 638 309 658 343
rect 544 283 658 309
rect 544 257 644 283
rect 104 81 204 107
rect 246 81 346 107
rect 402 81 502 107
rect 544 81 644 107
<< polycont >>
rect 110 317 144 351
rect 309 308 343 342
rect 425 309 459 343
rect 604 309 638 343
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 29 735 391 761
rect 29 701 45 735
rect 79 727 357 735
rect 79 701 95 727
rect 29 652 95 701
rect 341 701 357 727
rect 29 618 45 652
rect 79 618 95 652
rect 29 568 95 618
rect 29 534 45 568
rect 79 534 95 568
rect 29 485 95 534
rect 29 451 45 485
rect 79 451 95 485
rect 29 435 95 451
rect 185 657 201 691
rect 235 657 257 691
rect 185 623 257 657
rect 185 589 201 623
rect 235 589 257 623
rect 185 553 257 589
rect 185 519 201 553
rect 235 519 257 553
rect 185 485 257 519
rect 185 451 201 485
rect 235 451 257 485
rect 185 435 257 451
rect 25 351 167 367
rect 25 317 110 351
rect 144 317 167 351
rect 25 301 167 317
rect 18 249 136 265
rect 18 215 59 249
rect 93 215 136 249
rect 18 149 136 215
rect 217 196 257 435
rect 341 652 391 701
rect 341 618 357 652
rect 341 568 391 618
rect 341 534 357 568
rect 341 485 391 534
rect 341 451 357 485
rect 427 735 617 751
rect 427 701 433 735
rect 467 701 505 735
rect 547 701 577 735
rect 611 701 617 735
rect 427 654 617 701
rect 427 620 513 654
rect 547 620 617 654
rect 427 571 617 620
rect 427 537 513 571
rect 547 537 617 571
rect 427 490 617 537
rect 427 456 513 490
rect 547 456 617 490
rect 653 735 719 751
rect 653 701 669 735
rect 703 701 719 735
rect 653 652 719 701
rect 653 618 669 652
rect 703 618 719 652
rect 653 568 719 618
rect 653 534 669 568
rect 703 534 719 568
rect 653 485 719 534
rect 341 420 391 451
rect 653 451 669 485
rect 703 451 719 485
rect 653 420 719 451
rect 341 386 719 420
rect 293 342 359 350
rect 293 308 309 342
rect 343 308 359 342
rect 293 301 359 308
rect 409 343 551 350
rect 409 309 425 343
rect 459 309 551 343
rect 409 301 551 309
rect 588 343 743 350
rect 588 309 604 343
rect 638 309 743 343
rect 588 301 743 309
rect 341 249 391 265
rect 341 215 357 249
rect 341 196 391 215
rect 217 162 391 196
rect 18 115 59 149
rect 93 115 136 149
rect 18 113 136 115
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 136 113
rect 341 149 391 162
rect 341 115 357 149
rect 341 99 391 115
rect 427 249 750 265
rect 427 215 655 249
rect 689 215 750 249
rect 427 149 750 215
rect 427 115 655 149
rect 689 115 750 149
rect 427 113 750 115
rect 18 73 136 79
rect 461 79 499 113
rect 533 79 571 113
rect 605 79 643 113
rect 677 79 715 113
rect 749 79 750 113
rect 427 73 750 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 433 701 467 735
rect 505 701 513 735
rect 513 701 539 735
rect 577 701 611 735
rect 24 79 58 113
rect 96 79 130 113
rect 427 79 461 113
rect 499 79 533 113
rect 571 79 605 113
rect 643 79 677 113
rect 715 79 749 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 433 735
rect 467 701 505 735
rect 539 701 577 735
rect 611 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 427 113
rect 461 79 499 113
rect 533 79 571 113
rect 605 79 643 113
rect 677 79 715 113
rect 749 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a22oi_1
flabel metal1 s 0 51 768 125 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 0 768 23 0 FreeSans 340 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 0 689 768 763 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 791 768 814 0 FreeSans 340 0 0 0 VPB
port 7 nsew power bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 612 257 646 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 768 814
string GDS_END 794382
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 783900
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
