/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5.spice