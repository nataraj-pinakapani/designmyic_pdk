magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 3 11 4 6 DRAIN
port 1 nsew
rlabel  s 2 4 10 5 6 GATE
port 2 nsew
rlabel  s 2 0 10 1 8 GATE
port 2 nsew
rlabel  s 0 1 11 2 6 SOURCE
port 3 nsew
rlabel  s 0 1 1 4 4 SUBSTRATE
port 4 nsew
rlabel  s 11 1 11 4 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 11 5
string LEFview TRUE
<< end >>
