/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/lef/sky130_fd_io/sky130_ef_io.lef