magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< metal4 >>
rect 0 13600 1000 18593
rect 0 12410 1000 13300
rect 0 11240 1000 12130
rect 0 10874 1000 10940
rect 0 10218 1000 10814
rect 0 9266 1000 9862
rect 0 9140 1000 9206
rect 0 6940 1000 7630
rect 0 5970 1000 6660
rect 0 4760 1000 5690
rect 0 3550 1000 4480
rect 0 2580 1000 3270
rect 0 0 1000 1090
<< obsm4 >>
rect 0 34750 1000 39593
rect 0 9922 1000 10158
<< metal5 >>
rect 0 34750 1000 39593
rect 0 13600 1000 18590
rect 0 12430 1000 13280
rect 0 11260 1000 12110
rect 0 9140 1000 10940
rect 0 6960 1000 7610
rect 0 5990 1000 6640
rect 0 4780 1000 5670
rect 0 3570 1000 4460
rect 0 2600 1000 3250
rect 0 20 1000 1070
<< labels >>
rlabel metal4 s 0 10218 1000 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 1000 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 0 9140 1000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10874 1000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9140 1000 9206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6960 1000 7610 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6940 1000 7630 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 2600 1000 3250 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2580 1000 3270 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 5990 1000 6640 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 0 5970 1000 6660 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 0 12430 1000 13280 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 12410 1000 13300 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 20 1000 1070 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 0 0 1000 1090 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 13600 1000 18590 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 13600 1000 18593 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3570 1000 4460 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 3550 1000 4480 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 4780 1000 5670 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 0 4760 1000 5690 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 34750 1000 39593 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 11260 1000 12110 6 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 0 11240 1000 12130 6 VSSIO_Q
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1000 39593
string LEFclass PAD AREAIO
string LEFview TRUE
string GDS_END 8154
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_ef_io__disconnect_vccd_slice_5um.gds
string GDS_START 170
<< end >>
