magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel 
 s 1 93 14 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 93 14 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 93 14 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 92 15 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 92 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 92 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 92 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 92 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 92 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 92 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 91 16 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 91 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 91 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 91 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 91 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 91 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 90 17 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 90 17 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 90 17 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 90 17 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 90 17 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 90 17 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 90 17 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 89 18 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 89 18 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 89 18 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 89 18 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 89 18 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 89 18 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 89 18 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 88 19 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 88 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 88 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 88 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 88 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 88 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 87 20 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 87 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 87 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 87 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 87 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 87 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 87 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 86 21 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 86 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 86 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 86 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 86 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 86 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 86 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 85 22 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 85 22 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 85 22 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 85 22 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 85 22 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 85 22 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 84 23 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 84 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 84 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 84 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 84 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 84 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 84 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 83 24 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 83 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 83 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 83 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 83 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 83 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 68 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 18 25 22 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 51 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 61 93 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 61 93 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 61 93 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 61 92 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 61 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 60 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 60 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 60 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 60 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 60 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 60 91 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 59 91 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 59 91 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 59 91 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 59 91 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 59 91 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 59 90 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 59 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 58 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 58 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 58 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 58 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 58 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 58 89 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 58 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 57 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 57 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 57 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 57 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 57 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 57 88 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 56 88 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 56 88 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 56 88 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 56 88 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 56 88 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 56 87 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 56 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 55 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 55 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 55 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 55 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 55 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 55 86 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 55 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 54 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 54 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 54 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 54 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 54 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 54 85 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 53 85 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 53 85 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 53 85 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 53 85 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 53 85 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 53 84 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 53 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 52 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 52 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 52 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 52 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 52 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 52 83 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 52 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 51 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 51 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 51 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 51 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 51 68 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 18 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 93 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 83 14 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 83 1 83 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 25 83 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 68 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 14 91 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 14 88 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 14 83 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 16 88 18 90 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 19 86 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 19 83 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 22 83 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 93 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 68 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 61 83 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 51 68 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 51 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 52 83 54 84 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 54 83 56 86 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 55 86 56 87 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 56 83 61 88 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 58 88 59 90 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 59 88 61 91 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 60 91 61 92 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 22 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 22 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 21 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 21 75 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 75 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 75 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 75 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 19 75 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 19 75 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 18 75 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 18 75 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 93 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 92 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 75 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 75 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 90 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 75 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 75 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 88 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 88 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 75 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 75 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 86 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 85 75 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 85 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 75 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 75 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 83 75 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 82 74 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 82 74 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 82 74 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 81 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 81 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 80 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 80 74 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 80 74 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 79 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 79 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 78 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 78 74 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 78 74 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 77 74 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 77 74 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 76 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 76 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 75 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 75 74 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 75 74 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 74 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 74 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 73 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 73 74 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 73 74 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 72 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 72 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 71 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 71 74 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 71 74 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 70 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 70 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 69 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 69 74 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 69 74 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 68 74 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 22 74 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 22 74 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 21 74 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 21 74 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 74 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 74 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 74 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 19 74 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 19 74 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 93 74 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 92 74 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 92 74 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 74 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 74 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 74 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 90 74 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 90 74 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 74 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 74 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 74 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 88 74 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 88 74 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 74 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 74 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 74 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 86 74 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 86 74 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 85 74 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 85 74 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 74 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 74 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 74 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 83 74 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 83 74 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 82 74 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 82 74 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 82 74 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 81 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 81 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 80 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 80 74 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 80 74 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 79 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 79 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 78 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 78 74 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 78 74 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 77 74 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 77 74 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 76 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 76 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 75 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 75 74 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 75 74 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 74 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 74 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 73 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 73 74 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 73 74 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 72 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 72 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 71 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 71 74 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 71 74 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 70 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 70 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 69 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 69 74 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 69 74 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 68 74 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 22 74 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 22 74 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 21 74 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 21 74 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 74 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 74 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 20 74 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 19 74 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 19 74 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 18 74 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 93 74 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 92 74 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 92 74 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 74 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 74 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 91 74 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 90 74 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 90 74 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 74 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 74 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 89 74 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 88 74 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 88 74 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 74 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 74 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 87 74 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 86 74 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 86 74 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 85 74 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 85 74 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 74 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 74 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 84 74 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 83 74 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 74 83 74 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 74 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 74 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 74 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 81 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 81 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 74 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 74 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 74 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 79 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 79 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 74 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 74 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 74 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 77 74 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 77 74 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 76 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 76 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 74 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 74 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 74 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 74 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 74 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 74 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 74 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 74 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 72 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 72 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 74 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 74 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 74 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 70 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 70 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 74 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 74 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 74 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 68 74 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 22 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 22 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 21 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 21 73 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 20 73 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 20 73 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 20 73 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 19 73 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 19 73 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 93 73 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 92 73 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 92 73 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 91 73 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 91 73 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 91 73 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 90 73 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 90 73 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 89 73 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 89 73 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 89 73 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 88 73 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 88 73 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 87 73 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 87 73 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 87 73 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 86 73 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 86 73 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 85 73 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 85 73 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 84 73 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 84 73 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 84 73 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 83 73 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 83 73 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 73 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 73 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 73 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 81 73 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 81 73 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 73 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 73 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 73 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 79 73 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 79 73 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 73 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 73 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 73 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 77 73 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 77 73 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 76 73 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 76 73 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 73 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 73 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 73 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 74 73 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 74 73 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 73 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 73 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 73 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 72 73 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 72 73 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 73 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 73 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 73 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 70 73 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 70 73 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 73 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 73 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 73 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 68 73 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 22 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 22 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 21 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 21 73 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 20 73 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 20 73 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 20 73 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 19 73 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 19 73 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 18 73 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 93 73 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 92 73 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 92 73 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 91 73 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 91 73 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 91 73 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 90 73 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 90 73 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 89 73 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 89 73 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 89 73 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 88 73 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 88 73 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 87 73 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 87 73 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 87 73 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 86 73 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 86 73 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 85 73 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 85 73 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 84 73 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 84 73 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 84 73 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 83 73 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 83 73 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 73 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 73 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 82 73 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 81 73 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 81 73 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 73 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 73 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 80 73 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 79 73 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 79 73 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 73 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 73 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 78 73 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 77 73 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 77 73 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 76 73 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 76 73 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 73 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 73 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 75 73 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 74 73 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 74 73 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 73 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 73 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 73 73 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 72 73 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 72 73 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 73 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 73 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 71 73 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 70 73 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 70 73 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 73 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 73 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 69 73 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 73 68 73 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 22 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 22 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 21 73 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 21 73 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 73 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 73 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 73 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 19 73 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 19 73 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 18 73 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 18 73 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 93 72 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 92 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 92 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 91 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 91 72 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 91 72 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 90 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 90 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 89 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 89 72 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 89 72 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 88 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 88 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 87 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 87 72 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 87 72 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 86 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 86 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 85 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 85 72 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 84 72 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 84 72 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 84 72 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 83 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 83 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 82 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 82 72 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 82 72 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 81 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 81 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 80 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 80 72 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 80 72 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 79 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 79 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 78 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 78 72 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 78 72 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 77 72 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 77 72 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 76 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 76 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 75 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 75 72 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 75 72 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 74 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 74 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 73 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 73 72 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 73 72 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 72 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 72 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 71 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 71 72 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 71 72 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 70 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 70 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 69 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 69 72 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 69 72 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 68 72 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 22 72 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 22 72 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 21 72 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 21 72 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 72 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 72 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 72 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 19 72 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 19 72 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 93 72 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 92 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 92 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 91 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 91 72 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 91 72 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 90 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 90 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 89 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 89 72 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 89 72 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 88 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 88 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 87 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 87 72 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 87 72 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 86 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 86 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 85 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 85 72 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 84 72 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 84 72 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 84 72 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 83 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 83 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 82 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 82 72 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 82 72 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 81 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 81 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 80 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 80 72 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 80 72 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 79 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 79 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 78 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 78 72 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 78 72 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 77 72 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 77 72 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 76 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 76 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 75 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 75 72 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 75 72 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 74 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 74 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 73 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 73 72 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 73 72 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 72 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 72 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 71 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 71 72 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 71 72 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 70 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 70 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 69 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 69 72 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 69 72 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 68 72 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 22 72 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 22 72 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 21 72 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 21 72 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 72 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 72 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 20 72 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 19 72 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 19 72 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 72 18 72 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 93 72 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 92 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 92 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 72 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 72 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 72 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 90 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 90 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 72 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 72 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 72 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 88 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 88 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 72 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 72 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 72 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 86 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 86 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 85 72 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 85 72 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 72 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 72 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 72 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 83 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 83 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 72 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 72 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 72 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 81 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 81 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 72 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 72 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 72 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 79 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 79 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 72 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 72 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 72 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 77 72 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 77 72 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 76 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 76 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 72 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 72 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 72 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 74 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 74 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 72 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 72 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 72 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 72 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 72 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 72 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 72 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 72 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 70 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 70 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 72 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 72 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 72 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 68 72 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 22 71 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 22 71 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 21 71 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 21 71 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 20 71 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 20 71 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 20 71 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 19 71 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 19 71 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 93 71 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 92 71 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 92 71 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 71 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 71 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 71 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 90 71 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 90 71 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 71 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 71 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 71 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 88 71 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 88 71 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 71 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 71 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 71 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 86 71 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 86 71 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 85 71 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 85 71 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 71 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 71 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 71 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 83 71 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 83 71 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 71 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 71 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 71 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 81 71 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 81 71 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 71 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 71 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 71 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 79 71 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 79 71 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 71 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 71 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 71 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 77 71 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 77 71 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 76 71 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 76 71 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 71 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 71 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 71 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 74 71 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 74 71 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 71 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 71 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 71 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 72 71 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 72 71 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 71 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 71 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 71 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 70 71 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 70 71 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 71 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 71 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 71 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 68 71 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 22 71 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 22 71 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 21 71 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 21 71 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 20 71 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 20 71 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 20 71 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 19 71 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 19 71 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 18 71 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 93 71 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 92 71 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 92 71 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 71 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 71 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 91 71 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 90 71 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 90 71 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 71 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 71 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 89 71 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 88 71 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 88 71 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 71 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 71 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 87 71 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 86 71 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 86 71 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 85 71 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 85 71 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 71 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 71 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 84 71 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 83 71 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 83 71 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 71 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 71 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 82 71 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 81 71 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 81 71 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 71 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 71 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 80 71 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 79 71 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 79 71 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 71 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 71 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 78 71 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 77 71 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 77 71 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 76 71 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 76 71 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 71 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 71 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 75 71 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 74 71 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 74 71 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 71 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 71 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 73 71 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 72 71 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 72 71 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 71 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 71 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 71 71 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 70 71 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 70 71 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 71 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 71 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 69 71 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 71 68 71 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 22 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 22 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 21 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 21 70 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 20 70 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 20 70 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 20 70 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 19 70 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 19 70 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 93 70 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 92 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 92 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 91 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 91 70 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 91 70 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 90 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 90 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 89 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 89 70 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 89 70 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 88 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 88 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 87 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 87 70 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 87 70 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 86 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 86 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 85 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 85 70 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 84 70 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 84 70 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 84 70 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 83 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 83 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 82 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 82 70 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 82 70 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 81 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 81 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 80 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 80 70 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 80 70 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 79 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 79 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 78 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 78 70 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 78 70 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 77 70 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 77 70 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 76 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 76 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 75 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 75 70 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 75 70 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 74 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 74 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 73 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 73 70 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 73 70 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 72 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 72 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 71 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 71 70 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 71 70 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 70 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 70 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 69 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 69 70 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 69 70 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 68 70 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 22 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 22 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 21 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 21 70 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 20 70 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 20 70 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 20 70 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 19 70 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 19 70 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 18 70 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 93 70 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 92 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 92 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 91 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 91 70 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 91 70 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 90 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 90 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 89 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 89 70 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 89 70 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 88 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 88 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 87 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 87 70 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 87 70 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 86 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 86 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 85 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 85 70 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 84 70 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 84 70 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 84 70 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 83 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 83 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 82 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 82 70 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 82 70 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 81 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 81 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 80 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 80 70 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 80 70 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 79 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 79 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 78 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 78 70 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 78 70 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 77 70 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 77 70 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 76 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 76 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 75 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 75 70 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 75 70 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 74 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 74 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 73 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 73 70 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 73 70 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 72 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 72 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 71 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 71 70 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 71 70 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 70 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 70 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 69 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 69 70 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 69 70 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 70 68 70 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 22 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 22 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 21 70 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 21 70 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 70 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 70 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 70 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 19 70 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 19 70 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 18 70 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 18 70 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 70 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 70 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 81 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 81 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 70 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 70 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 70 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 79 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 79 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 70 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 70 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 70 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 77 70 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 77 70 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 76 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 76 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 70 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 70 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 70 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 74 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 74 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 70 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 70 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 70 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 72 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 72 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 70 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 70 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 70 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 70 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 70 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 70 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 70 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 70 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 68 70 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 93 70 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 92 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 92 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 70 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 70 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 70 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 90 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 90 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 70 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 70 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 70 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 88 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 88 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 70 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 70 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 70 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 86 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 86 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 85 70 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 85 70 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 70 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 70 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 70 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 83 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 83 70 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 22 69 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 22 69 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 21 69 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 21 69 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 69 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 69 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 69 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 19 69 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 19 69 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 69 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 69 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 69 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 81 69 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 81 69 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 69 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 69 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 69 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 79 69 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 79 69 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 69 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 69 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 69 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 77 69 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 77 69 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 76 69 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 76 69 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 69 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 69 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 69 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 74 69 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 74 69 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 69 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 69 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 69 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 72 69 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 72 69 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 69 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 69 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 69 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 70 69 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 70 69 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 69 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 69 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 69 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 68 69 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 93 69 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 92 69 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 92 69 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 69 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 69 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 69 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 90 69 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 90 69 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 69 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 69 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 69 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 88 69 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 88 69 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 69 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 69 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 69 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 86 69 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 86 69 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 85 69 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 85 69 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 69 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 69 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 69 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 83 69 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 83 69 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 22 69 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 22 69 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 21 69 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 21 69 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 69 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 69 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 20 69 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 19 69 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 19 69 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 18 69 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 69 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 69 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 82 69 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 81 69 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 81 69 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 69 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 69 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 80 69 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 79 69 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 79 69 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 69 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 69 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 78 69 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 77 69 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 77 69 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 76 69 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 76 69 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 69 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 69 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 75 69 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 74 69 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 74 69 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 69 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 69 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 73 69 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 72 69 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 72 69 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 69 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 69 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 71 69 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 70 69 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 70 69 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 69 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 69 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 69 69 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 68 69 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 93 69 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 92 69 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 92 69 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 69 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 69 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 91 69 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 90 69 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 90 69 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 69 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 69 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 89 69 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 88 69 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 88 69 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 69 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 69 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 87 69 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 86 69 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 86 69 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 85 69 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 85 69 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 69 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 69 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 84 69 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 83 69 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 69 83 69 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 22 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 22 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 21 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 21 68 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 20 68 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 20 68 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 20 68 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 19 68 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 19 68 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 82 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 82 68 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 82 68 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 81 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 81 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 80 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 80 68 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 80 68 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 79 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 79 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 78 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 78 68 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 78 68 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 77 68 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 77 68 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 76 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 76 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 75 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 75 68 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 75 68 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 74 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 74 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 73 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 73 68 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 73 68 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 72 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 72 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 71 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 71 68 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 71 68 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 70 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 70 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 69 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 69 68 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 69 68 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 68 68 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 93 68 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 92 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 92 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 91 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 91 68 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 91 68 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 90 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 90 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 89 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 89 68 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 89 68 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 88 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 88 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 87 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 87 68 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 87 68 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 86 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 86 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 85 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 85 68 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 84 68 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 84 68 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 84 68 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 83 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 83 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 22 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 22 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 21 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 21 68 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 20 68 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 20 68 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 20 68 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 19 68 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 19 68 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 18 68 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 82 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 82 68 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 82 68 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 81 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 81 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 80 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 80 68 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 80 68 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 79 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 79 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 78 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 78 68 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 78 68 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 77 68 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 77 68 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 76 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 76 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 75 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 75 68 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 75 68 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 74 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 74 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 73 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 73 68 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 73 68 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 72 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 72 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 71 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 71 68 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 71 68 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 70 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 70 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 69 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 69 68 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 69 68 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 68 68 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 93 68 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 92 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 92 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 91 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 91 68 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 91 68 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 90 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 90 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 89 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 89 68 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 89 68 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 88 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 88 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 87 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 87 68 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 87 68 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 86 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 86 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 85 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 85 68 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 84 68 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 84 68 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 84 68 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 83 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 68 83 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 22 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 22 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 21 68 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 21 68 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 68 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 68 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 68 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 19 68 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 19 68 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 18 68 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 18 68 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 68 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 68 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 81 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 81 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 68 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 68 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 68 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 79 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 79 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 68 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 68 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 68 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 77 68 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 77 68 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 76 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 76 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 68 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 68 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 68 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 74 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 74 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 68 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 68 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 68 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 72 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 72 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 68 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 68 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 68 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 70 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 70 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 68 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 68 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 68 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 68 68 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 93 68 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 92 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 92 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 68 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 68 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 68 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 90 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 90 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 68 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 68 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 68 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 88 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 88 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 68 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 68 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 68 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 86 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 86 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 85 68 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 85 68 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 68 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 68 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 68 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 83 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 83 68 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 22 67 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 22 67 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 21 67 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 21 67 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 67 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 67 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 67 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 19 67 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 19 67 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 67 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 67 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 67 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 81 67 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 81 67 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 67 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 67 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 67 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 79 67 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 79 67 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 67 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 67 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 67 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 77 67 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 77 67 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 76 67 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 76 67 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 67 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 67 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 67 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 74 67 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 74 67 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 67 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 67 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 67 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 72 67 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 72 67 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 67 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 67 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 67 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 70 67 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 70 67 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 67 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 67 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 67 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 68 67 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 93 67 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 92 67 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 92 67 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 67 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 67 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 67 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 90 67 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 90 67 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 67 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 67 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 67 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 88 67 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 88 67 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 67 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 67 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 67 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 86 67 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 86 67 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 85 67 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 85 67 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 67 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 67 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 67 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 83 67 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 83 67 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 22 67 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 22 67 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 21 67 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 21 67 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 67 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 67 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 20 67 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 19 67 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 19 67 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 18 67 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 67 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 67 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 82 67 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 81 67 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 81 67 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 67 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 67 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 80 67 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 79 67 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 79 67 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 67 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 67 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 78 67 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 77 67 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 77 67 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 76 67 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 76 67 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 67 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 67 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 75 67 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 74 67 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 74 67 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 67 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 67 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 73 67 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 72 67 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 72 67 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 67 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 67 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 71 67 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 70 67 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 70 67 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 67 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 67 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 69 67 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 68 67 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 93 67 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 92 67 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 92 67 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 67 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 67 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 91 67 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 90 67 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 90 67 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 67 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 67 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 89 67 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 88 67 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 88 67 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 67 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 67 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 87 67 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 86 67 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 86 67 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 85 67 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 85 67 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 67 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 67 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 84 67 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 83 67 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 67 83 67 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 22 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 22 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 21 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 21 66 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 20 66 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 20 66 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 20 66 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 19 66 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 19 66 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 18 66 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 18 66 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 82 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 82 66 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 82 66 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 81 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 81 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 80 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 80 66 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 80 66 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 79 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 79 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 78 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 78 66 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 78 66 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 77 66 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 77 66 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 76 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 76 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 75 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 75 66 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 75 66 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 74 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 74 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 73 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 73 66 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 73 66 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 72 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 72 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 71 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 71 66 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 71 66 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 70 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 70 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 69 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 69 66 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 69 66 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 68 66 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 93 66 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 92 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 92 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 91 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 91 66 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 91 66 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 90 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 90 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 89 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 89 66 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 89 66 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 88 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 88 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 87 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 87 66 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 87 66 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 86 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 86 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 85 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 85 66 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 84 66 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 84 66 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 84 66 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 83 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 83 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 22 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 22 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 21 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 21 66 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 20 66 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 20 66 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 20 66 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 19 66 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 19 66 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 18 66 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 18 66 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 82 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 82 66 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 82 66 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 81 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 81 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 80 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 80 66 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 80 66 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 79 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 79 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 78 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 78 66 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 78 66 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 77 66 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 77 66 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 76 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 76 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 75 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 75 66 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 75 66 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 74 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 74 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 73 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 73 66 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 73 66 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 72 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 72 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 71 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 71 66 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 71 66 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 70 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 70 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 69 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 69 66 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 69 66 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 68 66 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 93 66 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 92 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 92 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 91 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 91 66 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 91 66 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 90 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 90 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 89 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 89 66 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 89 66 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 88 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 88 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 87 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 87 66 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 87 66 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 86 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 86 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 85 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 85 66 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 84 66 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 84 66 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 84 66 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 83 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 66 83 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 22 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 22 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 21 66 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 21 66 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 66 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 66 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 66 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 19 66 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 19 66 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 18 66 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 18 66 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 66 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 66 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 81 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 81 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 66 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 66 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 66 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 79 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 79 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 66 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 66 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 66 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 77 66 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 77 66 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 76 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 76 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 66 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 66 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 66 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 74 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 74 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 66 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 66 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 66 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 72 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 72 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 66 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 66 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 66 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 70 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 70 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 66 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 66 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 66 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 68 66 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 93 66 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 92 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 92 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 91 66 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 91 66 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 91 66 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 90 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 90 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 89 66 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 89 66 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 89 66 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 88 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 88 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 87 66 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 87 66 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 87 66 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 86 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 86 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 85 66 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 85 66 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 84 66 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 84 66 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 84 66 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 83 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 83 66 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 22 65 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 22 65 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 21 65 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 21 65 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 65 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 65 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 65 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 19 65 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 19 65 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 65 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 65 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 65 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 81 65 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 81 65 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 65 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 65 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 65 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 79 65 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 79 65 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 65 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 65 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 65 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 77 65 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 77 65 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 76 65 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 76 65 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 65 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 65 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 65 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 74 65 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 74 65 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 65 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 65 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 65 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 72 65 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 72 65 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 65 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 65 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 65 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 70 65 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 70 65 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 65 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 65 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 65 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 68 65 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 93 65 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 92 65 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 92 65 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 91 65 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 91 65 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 91 65 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 90 65 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 90 65 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 89 65 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 89 65 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 89 65 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 88 65 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 88 65 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 87 65 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 87 65 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 87 65 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 86 65 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 86 65 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 85 65 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 85 65 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 84 65 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 84 65 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 84 65 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 83 65 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 83 65 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 22 65 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 22 65 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 21 65 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 21 65 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 65 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 65 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 20 65 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 19 65 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 19 65 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 18 65 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 65 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 65 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 82 65 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 81 65 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 81 65 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 65 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 65 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 80 65 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 79 65 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 79 65 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 65 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 65 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 78 65 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 77 65 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 77 65 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 76 65 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 76 65 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 65 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 65 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 75 65 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 74 65 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 74 65 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 65 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 65 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 73 65 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 72 65 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 72 65 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 65 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 65 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 71 65 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 70 65 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 70 65 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 65 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 65 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 69 65 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 65 68 65 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 93 65 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 92 65 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 92 65 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 65 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 65 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 65 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 90 65 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 90 65 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 65 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 65 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 65 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 88 65 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 88 65 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 65 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 65 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 65 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 86 65 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 86 65 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 85 65 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 85 65 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 65 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 65 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 65 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 83 65 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 83 65 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 82 64 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 82 64 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 82 64 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 81 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 81 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 80 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 80 64 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 80 64 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 79 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 79 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 78 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 78 64 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 78 64 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 77 64 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 77 64 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 76 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 76 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 75 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 75 64 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 75 64 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 74 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 74 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 73 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 73 64 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 73 64 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 72 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 72 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 71 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 71 64 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 71 64 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 70 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 70 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 69 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 69 64 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 69 64 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 68 64 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 22 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 22 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 21 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 21 64 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 20 64 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 20 64 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 20 64 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 19 64 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 19 64 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 93 64 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 92 64 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 92 64 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 64 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 64 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 64 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 90 64 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 90 64 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 64 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 64 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 64 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 88 64 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 88 64 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 64 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 64 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 64 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 86 64 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 86 64 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 85 64 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 85 64 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 64 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 64 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 64 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 83 64 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 83 64 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 82 64 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 82 64 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 82 64 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 81 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 81 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 80 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 80 64 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 80 64 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 79 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 79 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 78 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 78 64 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 78 64 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 77 64 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 77 64 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 76 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 76 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 75 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 75 64 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 75 64 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 74 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 74 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 73 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 73 64 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 73 64 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 72 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 72 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 71 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 71 64 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 71 64 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 70 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 70 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 69 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 69 64 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 69 64 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 68 64 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 22 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 22 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 21 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 21 64 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 20 64 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 20 64 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 20 64 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 19 64 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 19 64 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 18 64 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 93 64 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 92 64 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 92 64 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 64 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 64 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 91 64 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 90 64 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 90 64 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 64 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 64 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 89 64 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 88 64 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 88 64 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 64 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 64 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 87 64 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 86 64 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 86 64 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 85 64 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 85 64 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 64 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 64 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 84 64 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 83 64 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 64 83 64 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 64 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 64 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 64 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 81 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 81 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 64 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 64 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 64 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 79 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 79 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 64 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 64 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 64 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 77 64 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 77 64 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 76 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 76 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 64 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 64 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 64 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 74 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 74 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 64 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 64 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 64 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 72 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 72 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 64 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 64 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 64 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 70 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 70 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 64 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 64 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 64 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 68 64 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 22 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 22 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 21 64 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 21 64 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 64 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 64 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 64 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 19 64 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 19 64 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 18 64 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 18 64 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 93 63 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 92 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 92 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 91 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 91 63 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 91 63 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 90 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 90 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 89 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 89 63 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 89 63 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 88 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 88 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 87 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 87 63 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 87 63 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 86 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 86 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 85 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 85 63 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 84 63 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 84 63 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 84 63 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 83 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 83 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 63 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 63 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 81 63 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 81 63 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 63 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 63 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 63 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 79 63 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 79 63 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 63 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 63 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 63 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 77 63 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 77 63 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 76 63 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 76 63 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 63 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 63 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 63 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 74 63 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 74 63 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 63 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 63 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 63 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 72 63 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 72 63 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 63 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 63 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 63 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 70 63 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 70 63 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 63 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 63 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 63 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 68 63 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 22 63 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 22 63 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 21 63 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 21 63 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 63 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 63 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 63 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 19 63 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 19 63 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 93 63 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 92 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 92 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 91 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 91 63 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 91 63 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 90 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 90 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 89 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 89 63 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 89 63 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 88 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 88 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 87 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 87 63 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 87 63 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 86 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 86 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 85 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 85 63 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 84 63 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 84 63 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 84 63 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 83 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 83 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 63 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 82 63 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 81 63 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 81 63 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 63 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 63 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 80 63 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 79 63 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 79 63 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 63 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 63 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 78 63 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 77 63 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 77 63 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 76 63 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 76 63 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 63 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 63 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 75 63 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 74 63 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 74 63 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 63 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 63 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 73 63 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 72 63 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 72 63 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 63 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 63 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 71 63 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 70 63 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 70 63 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 63 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 63 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 69 63 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 68 63 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 22 63 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 22 63 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 21 63 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 21 63 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 63 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 63 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 20 63 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 19 63 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 19 63 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 63 18 63 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 93 63 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 92 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 92 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 63 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 63 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 63 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 90 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 90 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 63 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 63 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 63 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 88 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 88 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 63 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 63 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 63 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 86 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 86 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 85 63 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 85 63 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 63 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 63 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 63 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 83 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 83 63 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 82 62 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 82 62 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 82 62 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 81 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 81 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 80 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 80 62 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 80 62 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 79 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 79 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 78 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 78 62 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 78 62 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 77 62 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 77 62 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 76 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 76 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 75 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 75 62 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 75 62 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 74 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 74 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 73 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 73 62 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 73 62 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 72 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 72 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 71 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 71 62 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 71 62 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 70 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 70 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 69 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 69 62 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 69 62 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 68 62 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 22 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 22 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 21 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 21 62 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 20 62 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 20 62 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 20 62 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 19 62 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 19 62 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 93 62 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 92 62 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 92 62 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 62 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 62 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 62 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 90 62 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 90 62 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 62 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 62 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 62 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 88 62 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 88 62 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 62 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 62 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 62 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 86 62 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 86 62 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 85 62 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 85 62 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 62 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 62 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 62 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 83 62 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 83 62 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 82 62 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 82 62 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 82 62 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 81 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 81 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 80 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 80 62 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 80 62 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 79 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 79 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 78 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 78 62 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 78 62 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 77 62 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 77 62 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 76 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 76 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 75 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 75 62 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 75 62 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 74 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 74 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 73 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 73 62 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 73 62 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 72 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 72 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 71 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 71 62 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 71 62 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 70 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 70 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 69 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 69 62 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 69 62 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 68 62 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 22 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 22 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 21 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 21 62 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 20 62 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 20 62 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 20 62 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 19 62 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 19 62 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 18 62 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 93 62 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 92 62 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 92 62 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 62 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 62 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 91 62 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 90 62 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 90 62 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 62 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 62 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 89 62 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 88 62 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 88 62 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 62 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 62 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 87 62 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 86 62 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 86 62 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 85 62 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 85 62 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 62 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 62 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 84 62 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 83 62 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 62 83 62 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 62 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 62 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 62 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 81 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 81 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 62 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 62 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 62 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 79 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 79 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 62 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 62 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 62 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 77 62 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 77 62 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 76 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 76 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 62 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 62 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 62 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 74 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 74 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 62 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 62 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 62 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 72 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 72 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 62 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 62 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 62 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 70 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 70 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 62 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 62 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 62 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 68 62 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 22 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 22 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 21 62 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 21 62 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 62 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 62 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 62 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 19 62 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 19 62 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 18 62 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 18 62 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 93 61 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 92 61 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 92 61 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 91 61 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 91 61 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 91 61 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 90 61 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 90 61 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 89 61 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 89 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 89 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 88 61 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 88 61 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 87 61 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 87 61 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 87 61 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 86 61 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 86 61 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 85 61 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 85 61 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 84 61 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 84 61 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 84 61 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 83 61 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 83 61 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 61 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 61 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 61 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 81 61 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 81 61 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 61 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 61 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 61 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 79 61 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 79 61 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 61 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 61 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 61 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 77 61 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 77 61 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 76 61 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 76 61 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 61 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 61 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 61 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 74 61 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 74 61 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 61 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 61 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 61 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 72 61 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 72 61 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 61 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 61 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 61 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 70 61 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 70 61 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 61 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 61 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 61 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 68 61 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 22 61 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 22 61 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 21 61 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 21 61 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 61 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 61 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 61 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 19 61 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 19 61 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 91 61 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 91 61 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 91 61 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 90 61 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 90 61 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 89 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 89 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 88 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 61 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 61 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 82 61 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 81 61 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 81 61 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 61 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 61 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 80 61 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 79 61 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 79 61 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 61 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 61 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 78 61 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 77 61 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 77 61 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 76 61 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 76 61 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 61 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 61 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 75 61 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 74 61 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 74 61 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 61 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 61 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 73 61 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 72 61 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 72 61 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 61 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 61 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 71 61 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 70 61 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 70 61 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 61 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 61 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 69 61 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 68 61 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 88 61 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 87 61 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 87 61 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 87 61 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 86 61 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 86 61 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 85 61 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 85 61 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 85 61 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 84 61 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 84 61 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 83 61 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 83 61 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 22 61 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 22 61 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 21 61 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 21 61 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 61 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 61 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 20 61 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 19 61 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 19 61 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 61 18 61 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 91 61 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 90 61 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 90 61 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 89 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 89 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 88 61 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 82 60 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 82 60 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 82 60 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 81 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 81 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 80 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 80 60 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 80 60 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 79 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 79 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 78 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 78 60 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 78 60 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 77 60 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 77 60 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 76 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 76 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 75 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 75 60 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 75 60 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 74 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 74 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 73 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 73 60 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 73 60 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 72 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 72 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 71 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 71 60 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 71 60 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 70 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 70 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 69 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 69 60 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 69 60 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 68 60 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 88 60 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 87 60 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 87 60 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 87 60 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 86 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 86 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 85 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 85 60 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 85 60 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 84 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 84 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 83 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 83 60 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 22 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 22 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 21 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 21 60 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 20 60 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 20 60 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 20 60 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 19 60 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 19 60 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 91 60 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 91 60 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 91 60 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 90 60 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 90 60 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 89 60 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 89 60 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 88 60 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 82 60 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 82 60 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 82 60 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 81 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 81 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 80 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 80 60 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 80 60 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 79 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 79 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 78 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 78 60 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 78 60 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 77 60 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 77 60 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 76 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 76 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 75 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 75 60 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 75 60 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 74 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 74 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 73 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 73 60 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 73 60 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 72 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 72 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 71 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 71 60 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 71 60 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 70 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 70 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 69 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 69 60 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 69 60 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 68 60 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 88 60 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 87 60 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 87 60 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 87 60 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 86 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 86 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 85 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 85 60 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 85 60 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 84 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 84 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 83 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 83 60 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 22 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 22 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 21 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 21 60 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 20 60 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 20 60 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 20 60 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 19 60 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 19 60 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 60 18 60 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 91 60 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 90 60 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 90 60 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 89 60 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 89 60 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 88 60 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 60 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 60 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 60 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 81 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 81 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 60 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 60 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 60 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 79 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 79 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 60 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 60 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 60 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 77 60 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 77 60 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 76 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 76 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 60 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 60 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 60 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 74 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 74 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 60 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 60 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 60 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 72 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 72 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 60 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 60 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 60 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 70 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 70 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 60 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 60 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 60 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 68 60 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 88 60 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 60 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 60 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 60 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 86 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 86 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 60 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 60 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 60 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 84 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 84 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 83 60 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 83 60 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 22 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 22 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 21 60 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 21 60 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 60 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 60 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 60 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 19 60 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 19 60 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 18 60 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 18 60 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 91 59 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 90 59 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 90 59 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 89 59 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 89 59 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 88 59 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 59 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 59 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 59 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 81 59 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 81 59 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 59 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 59 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 59 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 79 59 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 79 59 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 59 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 59 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 59 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 77 59 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 77 59 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 76 59 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 76 59 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 59 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 59 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 59 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 74 59 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 74 59 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 59 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 59 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 59 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 72 59 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 72 59 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 59 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 59 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 59 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 70 59 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 70 59 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 59 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 59 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 59 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 68 59 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 88 59 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 59 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 59 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 59 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 86 59 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 86 59 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 59 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 59 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 59 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 84 59 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 84 59 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 83 59 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 83 59 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 22 59 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 22 59 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 21 59 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 21 59 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 59 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 59 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 59 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 19 59 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 19 59 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 59 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 59 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 82 59 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 81 59 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 81 59 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 59 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 59 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 80 59 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 79 59 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 79 59 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 59 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 59 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 78 59 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 77 59 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 77 59 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 76 59 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 76 59 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 59 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 59 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 75 59 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 74 59 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 74 59 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 59 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 59 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 73 59 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 72 59 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 72 59 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 59 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 59 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 71 59 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 70 59 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 70 59 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 59 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 59 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 69 59 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 68 59 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 89 59 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 89 59 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 88 59 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 88 59 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 59 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 59 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 87 59 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 86 59 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 86 59 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 59 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 59 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 85 59 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 84 59 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 84 59 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 83 59 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 83 59 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 22 59 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 22 59 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 21 59 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 21 59 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 59 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 59 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 20 59 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 19 59 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 19 59 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 59 18 59 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 82 58 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 82 58 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 82 58 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 81 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 81 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 80 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 80 58 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 80 58 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 79 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 79 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 78 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 78 58 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 78 58 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 77 58 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 77 58 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 76 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 76 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 75 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 75 58 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 75 58 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 74 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 74 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 73 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 73 58 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 73 58 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 72 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 72 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 71 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 71 58 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 71 58 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 70 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 70 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 69 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 69 58 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 69 58 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 68 58 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 22 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 22 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 21 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 21 58 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 20 58 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 20 58 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 20 58 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 19 58 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 19 58 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 88 58 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 87 58 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 87 58 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 87 58 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 86 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 86 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 85 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 85 58 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 85 58 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 84 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 84 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 83 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 83 58 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 82 58 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 82 58 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 82 58 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 81 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 81 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 80 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 80 58 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 80 58 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 79 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 79 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 78 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 78 58 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 78 58 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 77 58 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 77 58 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 76 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 76 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 75 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 75 58 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 75 58 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 74 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 74 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 73 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 73 58 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 73 58 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 72 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 72 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 71 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 71 58 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 71 58 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 70 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 70 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 69 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 69 58 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 69 58 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 68 58 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 89 58 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 89 58 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 88 58 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 22 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 22 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 21 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 21 58 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 20 58 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 20 58 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 20 58 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 19 58 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 19 58 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 18 58 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 88 58 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 87 58 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 87 58 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 87 58 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 86 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 86 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 85 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 85 58 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 85 58 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 84 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 84 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 83 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 58 83 58 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 58 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 58 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 58 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 81 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 81 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 58 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 58 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 58 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 79 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 79 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 58 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 58 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 58 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 77 58 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 77 58 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 76 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 76 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 58 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 58 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 58 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 74 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 74 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 58 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 58 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 58 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 72 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 72 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 58 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 58 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 58 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 70 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 70 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 58 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 58 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 58 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 68 58 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 22 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 22 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 21 58 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 21 58 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 58 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 58 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 58 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 19 58 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 19 58 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 18 58 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 18 58 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 88 58 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 87 58 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 87 58 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 87 58 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 86 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 86 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 85 58 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 85 58 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 85 58 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 84 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 84 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 83 58 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 83 58 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 57 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 57 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 57 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 81 57 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 81 57 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 57 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 57 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 57 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 79 57 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 79 57 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 57 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 57 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 57 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 77 57 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 77 57 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 76 57 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 76 57 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 57 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 57 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 57 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 74 57 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 74 57 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 57 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 57 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 57 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 72 57 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 72 57 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 57 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 57 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 57 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 70 57 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 70 57 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 57 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 57 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 57 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 68 57 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 22 57 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 22 57 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 21 57 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 21 57 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 57 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 57 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 57 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 19 57 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 19 57 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 88 57 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 87 57 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 87 57 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 87 57 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 86 57 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 86 57 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 85 57 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 85 57 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 85 57 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 84 57 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 84 57 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 83 57 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 83 57 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 57 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 57 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 82 57 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 81 57 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 81 57 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 57 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 57 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 80 57 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 79 57 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 79 57 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 57 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 57 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 78 57 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 77 57 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 77 57 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 76 57 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 76 57 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 57 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 57 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 75 57 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 74 57 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 74 57 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 57 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 57 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 73 57 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 72 57 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 72 57 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 57 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 57 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 71 57 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 70 57 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 70 57 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 57 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 57 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 69 57 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 68 57 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 22 57 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 22 57 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 21 57 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 21 57 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 57 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 57 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 20 57 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 19 57 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 19 57 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 57 18 57 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 88 57 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 87 57 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 87 57 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 87 57 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 86 57 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 86 57 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 85 57 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 85 57 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 85 57 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 84 57 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 84 57 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 83 57 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 83 57 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 82 56 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 82 56 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 82 56 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 81 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 81 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 80 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 80 56 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 80 56 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 79 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 79 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 78 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 78 56 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 78 56 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 77 56 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 77 56 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 76 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 76 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 75 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 75 56 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 75 56 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 74 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 74 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 73 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 73 56 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 73 56 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 72 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 72 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 71 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 71 56 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 71 56 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 70 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 70 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 69 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 69 56 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 69 56 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 68 56 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 22 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 22 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 21 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 21 56 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 20 56 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 20 56 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 20 56 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 19 56 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 19 56 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 87 56 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 86 56 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 86 56 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 82 56 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 82 56 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 82 56 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 81 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 81 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 80 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 80 56 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 80 56 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 79 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 79 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 78 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 78 56 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 78 56 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 77 56 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 77 56 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 76 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 76 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 75 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 75 56 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 75 56 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 74 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 74 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 73 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 73 56 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 73 56 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 72 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 72 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 71 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 71 56 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 71 56 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 70 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 70 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 69 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 69 56 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 69 56 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 68 56 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 85 56 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 85 56 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 84 56 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 84 56 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 83 56 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 83 56 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 22 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 22 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 21 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 21 56 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 20 56 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 20 56 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 20 56 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 19 56 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 19 56 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 56 18 56 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 56 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 56 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 56 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 81 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 81 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 56 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 56 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 56 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 79 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 79 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 56 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 56 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 56 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 77 56 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 77 56 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 76 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 76 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 56 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 56 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 56 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 74 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 74 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 56 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 56 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 56 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 72 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 72 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 56 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 56 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 56 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 70 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 70 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 56 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 56 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 56 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 68 56 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 85 56 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 85 56 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 84 56 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 84 56 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 83 56 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 83 56 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 22 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 22 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 21 56 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 21 56 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 20 56 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 20 56 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 20 56 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 19 56 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 19 56 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 18 56 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 18 56 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 87 55 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 86 55 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 86 55 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 55 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 55 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 55 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 81 55 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 81 55 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 55 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 55 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 55 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 79 55 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 79 55 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 55 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 55 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 55 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 77 55 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 77 55 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 76 55 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 76 55 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 55 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 55 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 55 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 74 55 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 74 55 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 55 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 55 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 55 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 72 55 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 72 55 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 55 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 55 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 55 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 70 55 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 70 55 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 55 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 55 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 55 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 68 55 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 22 55 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 22 55 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 21 55 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 21 55 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 20 55 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 20 55 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 20 55 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 19 55 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 19 55 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 18 55 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 18 55 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 85 55 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 85 55 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 84 55 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 84 55 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 83 55 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 83 55 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 55 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 55 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 82 55 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 81 55 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 81 55 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 55 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 55 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 80 55 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 79 55 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 79 55 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 55 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 55 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 78 55 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 77 55 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 77 55 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 76 55 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 76 55 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 55 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 55 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 75 55 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 74 55 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 74 55 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 55 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 55 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 73 55 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 72 55 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 72 55 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 55 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 55 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 71 55 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 70 55 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 70 55 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 55 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 55 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 69 55 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 55 68 55 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 22 55 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 22 55 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 21 55 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 21 55 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 55 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 55 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 55 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 19 55 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 19 55 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 18 55 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 18 55 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 85 55 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 85 55 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 84 55 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 84 55 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 83 55 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 83 55 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 82 54 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 82 54 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 82 54 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 81 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 81 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 80 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 80 54 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 80 54 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 79 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 79 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 78 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 78 54 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 78 54 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 77 54 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 77 54 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 76 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 76 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 75 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 75 54 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 75 54 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 74 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 74 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 73 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 73 54 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 73 54 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 72 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 72 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 71 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 71 54 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 71 54 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 70 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 70 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 69 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 69 54 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 69 54 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 68 54 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 22 54 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 22 54 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 21 54 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 21 54 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 54 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 54 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 54 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 19 54 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 19 54 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 85 54 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 85 54 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 84 54 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 84 54 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 83 54 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 83 54 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 82 54 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 82 54 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 82 54 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 81 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 81 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 80 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 80 54 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 80 54 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 79 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 79 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 78 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 78 54 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 78 54 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 77 54 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 77 54 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 76 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 76 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 75 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 75 54 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 75 54 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 74 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 74 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 73 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 73 54 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 73 54 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 72 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 72 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 71 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 71 54 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 71 54 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 70 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 70 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 69 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 69 54 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 69 54 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 68 54 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 22 54 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 22 54 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 21 54 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 21 54 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 54 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 54 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 20 54 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 19 54 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 19 54 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 54 18 54 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 54 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 54 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 54 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 81 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 81 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 54 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 54 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 54 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 79 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 79 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 54 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 54 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 54 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 77 54 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 77 54 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 76 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 76 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 54 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 54 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 54 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 74 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 74 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 54 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 54 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 54 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 72 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 72 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 54 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 54 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 54 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 70 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 70 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 54 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 54 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 54 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 68 54 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 84 54 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 83 54 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 83 54 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 22 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 22 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 21 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 21 53 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 20 53 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 20 53 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 20 53 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 19 53 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 19 53 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 53 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 53 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 53 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 81 53 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 81 53 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 53 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 53 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 53 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 79 53 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 79 53 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 53 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 53 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 53 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 77 53 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 77 53 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 76 53 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 76 53 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 53 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 53 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 53 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 74 53 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 74 53 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 53 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 53 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 53 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 72 53 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 72 53 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 53 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 53 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 53 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 70 53 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 70 53 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 53 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 53 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 53 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 68 53 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 22 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 22 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 21 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 21 53 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 20 53 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 20 53 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 20 53 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 19 53 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 19 53 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 18 53 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 53 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 53 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 82 53 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 81 53 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 81 53 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 53 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 53 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 80 53 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 79 53 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 79 53 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 53 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 53 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 78 53 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 77 53 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 77 53 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 76 53 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 76 53 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 53 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 53 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 75 53 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 74 53 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 74 53 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 53 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 53 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 73 53 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 72 53 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 72 53 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 53 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 53 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 71 53 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 70 53 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 70 53 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 53 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 53 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 69 53 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 68 53 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 84 53 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 83 53 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 53 83 53 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 22 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 22 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 21 53 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 21 53 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 53 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 53 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 53 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 19 53 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 19 53 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 18 53 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 18 53 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 82 52 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 82 52 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 82 52 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 81 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 81 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 80 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 80 52 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 80 52 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 79 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 79 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 78 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 78 52 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 78 52 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 77 52 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 77 52 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 76 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 76 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 75 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 75 52 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 75 52 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 74 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 74 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 73 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 73 52 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 73 52 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 72 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 72 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 71 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 71 52 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 71 52 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 70 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 70 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 69 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 69 52 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 69 52 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 68 52 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 22 52 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 22 52 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 21 52 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 21 52 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 52 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 52 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 52 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 19 52 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 19 52 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 82 52 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 82 52 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 82 52 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 81 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 81 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 80 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 80 52 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 80 52 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 79 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 79 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 78 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 78 52 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 78 52 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 77 52 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 77 52 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 76 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 76 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 75 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 75 52 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 75 52 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 74 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 74 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 73 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 73 52 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 73 52 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 72 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 72 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 71 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 71 52 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 71 52 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 70 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 70 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 69 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 69 52 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 69 52 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 68 52 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 22 52 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 22 52 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 21 52 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 21 52 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 52 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 52 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 20 52 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 19 52 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 19 52 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 52 18 52 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 82 52 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 82 52 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 82 52 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 81 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 81 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 80 52 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 80 52 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 80 52 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 79 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 79 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 78 52 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 78 52 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 78 52 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 77 52 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 77 52 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 76 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 76 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 75 52 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 75 52 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 75 52 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 74 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 74 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 73 52 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 73 52 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 73 52 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 72 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 72 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 71 52 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 71 52 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 71 52 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 70 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 70 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 69 52 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 69 52 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 69 52 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 68 52 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 22 51 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 22 51 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 21 51 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 21 51 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 20 51 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 20 51 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 20 51 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 19 51 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 19 51 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 18 51 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 18 51 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 82 51 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 82 51 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 82 51 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 81 51 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 81 51 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 80 51 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 80 51 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 80 51 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 79 51 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 79 51 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 78 51 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 78 51 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 78 51 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 77 51 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 77 51 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 76 51 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 76 51 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 75 51 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 75 51 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 75 51 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 74 51 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 74 51 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 73 51 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 73 51 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 73 51 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 72 51 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 72 51 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 71 51 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 71 51 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 71 51 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 70 51 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 70 51 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 69 51 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 69 51 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 69 51 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 68 51 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 22 51 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 22 51 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 21 51 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 21 51 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 20 51 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 20 51 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 20 51 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 19 51 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 19 51 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 18 51 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 51 18 51 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 22 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 22 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 21 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 21 24 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 20 24 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 20 24 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 20 24 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 19 24 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 19 24 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 82 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 82 24 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 82 24 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 81 24 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 81 24 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 80 24 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 80 24 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 80 24 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 79 24 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 79 24 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 78 24 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 78 24 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 78 24 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 77 24 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 77 24 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 76 24 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 76 24 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 75 24 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 75 24 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 75 24 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 74 24 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 74 24 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 73 24 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 73 24 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 73 24 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 72 24 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 72 24 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 71 24 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 71 24 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 71 24 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 70 24 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 70 24 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 69 24 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 69 24 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 69 24 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 68 24 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 22 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 22 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 21 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 21 24 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 20 24 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 20 24 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 20 24 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 19 24 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 19 24 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 18 24 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 82 24 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 82 24 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 82 24 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 81 24 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 81 24 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 80 24 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 80 24 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 80 24 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 79 24 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 79 24 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 78 24 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 78 24 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 78 24 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 77 24 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 77 24 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 76 24 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 76 24 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 75 24 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 75 24 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 75 24 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 74 24 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 74 24 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 73 24 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 73 24 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 73 24 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 72 24 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 72 24 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 71 24 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 71 24 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 71 24 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 70 24 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 70 24 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 69 24 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 69 24 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 69 24 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 24 68 24 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 22 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 22 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 21 24 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 21 24 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 24 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 24 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 24 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 19 24 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 19 24 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 18 24 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 18 24 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 82 23 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 82 23 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 82 23 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 81 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 81 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 80 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 80 23 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 80 23 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 79 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 79 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 78 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 78 23 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 78 23 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 77 23 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 77 23 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 76 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 76 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 75 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 75 23 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 75 23 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 74 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 74 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 73 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 73 23 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 73 23 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 72 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 72 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 71 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 71 23 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 71 23 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 70 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 70 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 69 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 69 23 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 69 23 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 68 23 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 22 23 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 22 23 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 21 23 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 21 23 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 23 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 23 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 23 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 19 23 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 19 23 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 82 23 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 82 23 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 82 23 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 81 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 81 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 80 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 80 23 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 80 23 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 79 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 79 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 78 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 78 23 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 78 23 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 77 23 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 77 23 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 76 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 76 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 75 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 75 23 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 75 23 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 74 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 74 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 73 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 73 23 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 73 23 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 72 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 72 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 71 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 71 23 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 71 23 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 70 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 70 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 69 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 69 23 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 69 23 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 68 23 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 22 23 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 22 23 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 21 23 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 21 23 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 23 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 23 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 20 23 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 19 23 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 19 23 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 18 23 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 84 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 83 23 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 23 83 23 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 23 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 23 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 23 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 81 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 81 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 23 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 23 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 23 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 79 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 79 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 23 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 23 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 23 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 77 23 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 77 23 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 76 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 76 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 23 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 23 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 23 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 74 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 74 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 23 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 23 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 23 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 72 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 72 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 23 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 23 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 23 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 70 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 70 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 23 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 23 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 23 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 68 23 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 22 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 22 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 21 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 21 22 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 20 22 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 20 22 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 20 22 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 19 22 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 19 22 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 22 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 22 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 22 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 81 22 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 81 22 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 22 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 22 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 22 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 79 22 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 79 22 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 22 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 22 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 22 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 77 22 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 77 22 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 76 22 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 76 22 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 22 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 22 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 22 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 74 22 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 74 22 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 22 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 22 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 22 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 72 22 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 72 22 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 22 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 22 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 22 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 70 22 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 70 22 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 22 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 22 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 22 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 68 22 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 22 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 22 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 21 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 21 22 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 20 22 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 20 22 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 20 22 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 19 22 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 19 22 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 18 22 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 84 22 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 83 22 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 83 22 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 22 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 22 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 82 22 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 81 22 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 81 22 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 22 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 22 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 80 22 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 79 22 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 79 22 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 22 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 22 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 78 22 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 77 22 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 77 22 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 76 22 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 76 22 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 22 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 22 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 75 22 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 74 22 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 74 22 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 22 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 22 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 73 22 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 72 22 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 72 22 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 22 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 22 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 71 22 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 70 22 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 70 22 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 22 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 22 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 69 22 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 22 68 22 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 22 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 22 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 21 22 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 21 22 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 22 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 22 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 22 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 19 22 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 19 22 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 18 22 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 18 22 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 82 21 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 82 21 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 82 21 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 81 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 81 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 80 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 80 21 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 80 21 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 79 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 79 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 78 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 78 21 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 78 21 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 77 21 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 77 21 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 76 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 76 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 75 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 75 21 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 75 21 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 74 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 74 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 73 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 73 21 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 73 21 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 72 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 72 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 71 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 71 21 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 71 21 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 70 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 70 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 69 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 69 21 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 69 21 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 68 21 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 85 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 85 21 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 84 21 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 84 21 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 83 21 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 83 21 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 22 21 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 22 21 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 21 21 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 21 21 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 21 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 21 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 21 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 19 21 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 19 21 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 82 21 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 82 21 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 82 21 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 81 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 81 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 80 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 80 21 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 80 21 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 79 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 79 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 78 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 78 21 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 78 21 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 77 21 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 77 21 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 76 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 76 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 75 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 75 21 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 75 21 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 74 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 74 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 73 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 73 21 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 73 21 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 72 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 72 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 71 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 71 21 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 71 21 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 70 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 70 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 69 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 69 21 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 69 21 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 68 21 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 85 21 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 85 21 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 84 21 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 84 21 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 83 21 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 83 21 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 22 21 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 22 21 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 21 21 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 21 21 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 21 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 21 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 20 21 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 19 21 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 19 21 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 21 18 21 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 21 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 21 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 21 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 81 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 81 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 21 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 21 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 21 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 79 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 79 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 21 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 21 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 21 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 77 21 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 77 21 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 76 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 76 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 21 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 21 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 21 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 74 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 74 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 21 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 21 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 21 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 72 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 72 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 21 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 21 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 21 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 70 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 70 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 21 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 21 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 21 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 68 21 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 85 20 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 85 20 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 84 20 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 84 20 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 83 20 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 83 20 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 22 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 22 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 21 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 21 20 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 20 20 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 20 20 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 20 20 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 19 20 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 19 20 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 20 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 20 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 20 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 81 20 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 81 20 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 20 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 20 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 20 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 79 20 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 79 20 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 20 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 20 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 20 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 77 20 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 77 20 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 76 20 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 76 20 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 20 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 20 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 20 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 74 20 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 74 20 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 20 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 20 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 20 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 72 20 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 72 20 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 20 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 20 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 20 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 70 20 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 70 20 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 20 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 20 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 20 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 68 20 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 87 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 86 20 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 86 20 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 85 20 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 85 20 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 84 20 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 84 20 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 83 20 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 83 20 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 22 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 22 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 21 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 21 20 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 20 20 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 20 20 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 20 20 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 19 20 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 19 20 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 18 20 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 20 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 20 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 82 20 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 81 20 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 81 20 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 20 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 20 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 80 20 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 79 20 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 79 20 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 20 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 20 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 78 20 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 77 20 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 77 20 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 76 20 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 76 20 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 20 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 20 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 75 20 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 74 20 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 74 20 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 20 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 20 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 73 20 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 72 20 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 72 20 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 20 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 20 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 71 20 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 70 20 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 70 20 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 20 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 20 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 69 20 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 20 68 20 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 22 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 22 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 21 20 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 21 20 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 20 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 20 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 20 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 19 20 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 19 20 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 18 20 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 18 20 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 85 19 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 85 19 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 84 19 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 84 19 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 83 19 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 83 19 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 82 19 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 82 19 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 82 19 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 81 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 81 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 80 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 80 19 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 80 19 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 79 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 79 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 78 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 78 19 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 78 19 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 77 19 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 77 19 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 76 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 76 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 75 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 75 19 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 75 19 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 74 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 74 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 73 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 73 19 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 73 19 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 72 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 72 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 71 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 71 19 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 71 19 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 70 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 70 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 69 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 69 19 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 69 19 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 68 19 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 87 19 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 86 19 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 86 19 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 22 19 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 22 19 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 21 19 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 21 19 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 19 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 19 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 19 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 19 19 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 19 19 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 82 19 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 82 19 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 82 19 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 81 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 81 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 80 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 80 19 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 80 19 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 79 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 79 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 78 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 78 19 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 78 19 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 77 19 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 77 19 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 76 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 76 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 75 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 75 19 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 75 19 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 74 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 74 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 73 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 73 19 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 73 19 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 72 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 72 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 71 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 71 19 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 71 19 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 70 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 70 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 69 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 69 19 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 69 19 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 68 19 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 88 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 87 19 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 87 19 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 87 19 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 86 19 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 86 19 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 85 19 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 85 19 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 85 19 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 84 19 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 84 19 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 83 19 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 83 19 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 22 19 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 22 19 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 21 19 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 21 19 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 19 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 19 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 20 19 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 19 19 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 19 19 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 19 18 19 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 19 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 19 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 19 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 81 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 81 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 19 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 19 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 19 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 79 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 79 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 19 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 19 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 19 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 77 19 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 77 19 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 76 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 76 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 19 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 19 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 19 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 74 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 74 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 19 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 19 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 19 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 72 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 72 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 19 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 19 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 19 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 70 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 70 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 19 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 19 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 19 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 68 19 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 88 18 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 87 18 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 87 18 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 87 18 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 86 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 86 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 85 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 85 18 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 85 18 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 84 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 84 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 83 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 83 18 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 22 18 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 22 18 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 21 18 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 21 18 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 20 18 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 20 18 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 20 18 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 19 18 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 19 18 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 18 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 18 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 18 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 81 18 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 81 18 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 18 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 18 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 18 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 79 18 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 79 18 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 18 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 18 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 18 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 77 18 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 77 18 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 76 18 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 76 18 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 18 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 18 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 18 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 74 18 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 74 18 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 18 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 18 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 18 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 72 18 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 72 18 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 18 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 18 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 18 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 70 18 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 70 18 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 18 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 18 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 18 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 68 18 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 88 18 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 87 18 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 87 18 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 87 18 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 86 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 86 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 85 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 85 18 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 85 18 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 84 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 84 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 83 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 83 18 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 22 18 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 22 18 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 21 18 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 21 18 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 20 18 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 20 18 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 20 18 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 19 18 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 19 18 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 18 18 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 18 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 18 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 82 18 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 81 18 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 81 18 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 18 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 18 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 80 18 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 79 18 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 79 18 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 18 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 18 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 78 18 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 77 18 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 77 18 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 76 18 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 76 18 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 18 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 18 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 75 18 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 74 18 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 74 18 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 18 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 18 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 73 18 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 72 18 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 72 18 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 18 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 18 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 71 18 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 70 18 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 70 18 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 18 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 18 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 69 18 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 18 68 18 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 88 18 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 18 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 18 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 18 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 86 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 86 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 18 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 18 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 18 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 84 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 84 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 83 18 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 83 18 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 22 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 22 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 21 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 21 17 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 20 17 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 20 17 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 20 17 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 19 17 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 19 17 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 89 17 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 89 17 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 88 17 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 82 17 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 82 17 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 82 17 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 81 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 81 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 80 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 80 17 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 80 17 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 79 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 79 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 78 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 78 17 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 78 17 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 77 17 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 77 17 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 76 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 76 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 75 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 75 17 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 75 17 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 74 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 74 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 73 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 73 17 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 73 17 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 72 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 72 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 71 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 71 17 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 71 17 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 70 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 70 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 69 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 69 17 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 69 17 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 68 17 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 88 17 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 17 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 17 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 17 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 86 17 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 86 17 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 17 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 17 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 17 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 84 17 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 84 17 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 83 17 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 83 17 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 22 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 22 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 21 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 21 17 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 20 17 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 20 17 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 20 17 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 19 17 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 19 17 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 18 17 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 82 17 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 82 17 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 82 17 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 81 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 81 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 80 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 80 17 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 80 17 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 79 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 79 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 78 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 78 17 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 78 17 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 77 17 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 77 17 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 76 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 76 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 75 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 75 17 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 75 17 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 74 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 74 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 73 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 73 17 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 73 17 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 72 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 72 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 71 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 71 17 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 71 17 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 70 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 70 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 69 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 69 17 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 69 17 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 68 17 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 88 17 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 17 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 17 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 87 17 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 86 17 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 86 17 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 17 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 17 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 85 17 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 84 17 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 84 17 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 83 17 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 17 83 17 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 22 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 22 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 21 17 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 21 17 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 17 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 17 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 17 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 19 17 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 19 17 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 18 17 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 18 17 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 89 17 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 89 17 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 88 17 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 17 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 17 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 17 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 81 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 81 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 17 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 17 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 17 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 79 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 79 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 17 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 17 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 17 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 77 17 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 77 17 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 76 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 76 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 17 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 17 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 17 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 74 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 74 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 17 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 17 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 17 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 72 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 72 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 17 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 17 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 17 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 70 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 70 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 17 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 17 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 17 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 68 17 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 88 16 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 87 16 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 87 16 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 87 16 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 86 16 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 86 16 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 85 16 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 85 16 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 85 16 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 84 16 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 84 16 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 83 16 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 83 16 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 22 16 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 22 16 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 21 16 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 21 16 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 16 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 16 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 16 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 19 16 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 19 16 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 16 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 16 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 16 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 81 16 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 81 16 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 16 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 16 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 16 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 79 16 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 79 16 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 16 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 16 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 16 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 77 16 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 77 16 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 76 16 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 76 16 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 16 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 16 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 16 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 74 16 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 74 16 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 16 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 16 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 16 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 72 16 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 72 16 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 16 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 16 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 16 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 70 16 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 70 16 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 16 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 16 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 16 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 68 16 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 91 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 90 16 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 90 16 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 89 16 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 89 16 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 88 16 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 88 16 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 87 16 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 87 16 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 87 16 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 86 16 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 86 16 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 85 16 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 85 16 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 85 16 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 84 16 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 84 16 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 83 16 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 83 16 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 22 16 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 22 16 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 21 16 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 21 16 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 16 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 16 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 20 16 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 19 16 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 19 16 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 18 16 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 16 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 16 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 82 16 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 81 16 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 81 16 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 16 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 16 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 80 16 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 79 16 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 79 16 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 16 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 16 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 78 16 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 77 16 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 77 16 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 76 16 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 76 16 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 16 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 16 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 75 16 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 74 16 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 74 16 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 16 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 16 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 73 16 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 72 16 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 72 16 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 16 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 16 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 71 16 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 70 16 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 70 16 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 16 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 16 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 69 16 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 68 16 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 91 16 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 90 16 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 90 16 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 89 16 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 89 16 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 16 88 16 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 88 15 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 87 15 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 87 15 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 87 15 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 86 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 86 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 85 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 85 15 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 85 15 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 84 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 84 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 83 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 83 15 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 22 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 22 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 21 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 21 15 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 20 15 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 20 15 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 20 15 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 19 15 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 19 15 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 82 15 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 82 15 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 82 15 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 81 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 81 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 80 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 80 15 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 80 15 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 79 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 79 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 78 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 78 15 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 78 15 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 77 15 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 77 15 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 76 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 76 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 75 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 75 15 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 75 15 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 74 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 74 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 73 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 73 15 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 73 15 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 72 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 72 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 71 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 71 15 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 71 15 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 70 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 70 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 69 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 69 15 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 69 15 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 68 15 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 91 15 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 90 15 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 90 15 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 89 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 89 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 88 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 91 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 91 15 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 88 15 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 87 15 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 87 15 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 87 15 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 86 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 86 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 85 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 85 15 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 85 15 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 84 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 84 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 83 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 83 15 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 22 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 22 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 21 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 21 15 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 20 15 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 20 15 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 20 15 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 19 15 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 19 15 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 18 15 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 82 15 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 82 15 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 82 15 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 81 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 81 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 80 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 80 15 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 80 15 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 79 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 79 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 78 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 78 15 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 78 15 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 77 15 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 77 15 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 76 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 76 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 75 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 75 15 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 75 15 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 74 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 74 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 73 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 73 15 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 73 15 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 72 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 72 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 71 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 71 15 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 71 15 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 70 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 70 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 69 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 69 15 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 69 15 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 68 15 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 91 15 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 90 15 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 90 15 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 89 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 89 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 15 88 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 88 15 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 87 15 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 87 15 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 87 15 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 86 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 86 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 85 15 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 85 15 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 85 15 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 84 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 84 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 83 15 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 83 15 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 22 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 22 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 21 15 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 21 15 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 15 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 15 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 15 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 19 15 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 19 15 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 18 15 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 18 15 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 15 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 15 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 15 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 81 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 81 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 15 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 15 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 15 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 79 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 79 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 15 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 15 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 15 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 77 15 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 77 15 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 76 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 76 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 15 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 15 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 15 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 74 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 74 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 15 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 15 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 15 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 72 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 72 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 15 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 15 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 15 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 70 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 70 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 15 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 15 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 15 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 68 15 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 91 15 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 90 15 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 90 15 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 89 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 89 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 88 15 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 91 15 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 91 15 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 22 14 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 22 14 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 21 14 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 21 14 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 14 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 14 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 14 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 19 14 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 19 14 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 14 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 14 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 14 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 81 14 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 81 14 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 14 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 14 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 14 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 79 14 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 79 14 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 14 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 14 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 14 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 77 14 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 77 14 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 76 14 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 76 14 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 14 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 14 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 14 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 74 14 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 74 14 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 14 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 14 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 14 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 72 14 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 72 14 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 14 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 14 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 14 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 70 14 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 70 14 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 14 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 14 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 14 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 68 14 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 93 14 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 92 14 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 92 14 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 91 14 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 91 14 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 91 14 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 90 14 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 90 14 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 89 14 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 89 14 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 89 14 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 88 14 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 88 14 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 87 14 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 87 14 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 87 14 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 86 14 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 86 14 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 85 14 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 85 14 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 84 14 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 84 14 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 84 14 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 83 14 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 83 14 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 22 14 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 22 14 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 21 14 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 21 14 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 14 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 14 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 20 14 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 19 14 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 19 14 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 18 14 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 14 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 14 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 82 14 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 81 14 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 81 14 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 14 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 14 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 80 14 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 79 14 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 79 14 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 14 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 14 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 78 14 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 77 14 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 77 14 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 76 14 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 76 14 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 14 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 14 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 75 14 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 74 14 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 74 14 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 14 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 14 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 73 14 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 72 14 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 72 14 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 14 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 14 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 71 14 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 70 14 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 70 14 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 14 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 14 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 69 14 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 14 68 14 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 93 14 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 92 14 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 92 14 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 14 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 14 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 14 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 90 14 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 90 14 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 14 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 14 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 14 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 88 14 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 88 14 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 14 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 14 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 14 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 86 14 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 86 14 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 85 14 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 85 14 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 14 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 14 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 14 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 83 14 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 83 14 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 82 13 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 82 13 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 82 13 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 81 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 81 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 80 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 80 13 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 80 13 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 79 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 79 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 78 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 78 13 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 78 13 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 77 13 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 77 13 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 76 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 76 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 75 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 75 13 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 75 13 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 74 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 74 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 73 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 73 13 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 73 13 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 72 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 72 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 71 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 71 13 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 71 13 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 70 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 70 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 69 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 69 13 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 69 13 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 68 13 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 22 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 22 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 21 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 21 13 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 20 13 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 20 13 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 20 13 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 19 13 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 19 13 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 93 13 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 92 13 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 92 13 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 13 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 13 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 13 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 90 13 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 90 13 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 13 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 13 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 13 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 88 13 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 88 13 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 13 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 13 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 13 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 86 13 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 86 13 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 85 13 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 85 13 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 13 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 13 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 13 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 83 13 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 83 13 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 82 13 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 82 13 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 82 13 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 81 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 81 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 80 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 80 13 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 80 13 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 79 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 79 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 78 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 78 13 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 78 13 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 77 13 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 77 13 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 76 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 76 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 75 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 75 13 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 75 13 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 74 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 74 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 73 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 73 13 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 73 13 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 72 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 72 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 71 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 71 13 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 71 13 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 70 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 70 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 69 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 69 13 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 69 13 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 68 13 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 22 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 22 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 21 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 21 13 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 20 13 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 20 13 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 20 13 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 19 13 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 19 13 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 18 13 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 93 13 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 92 13 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 92 13 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 13 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 13 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 91 13 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 90 13 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 90 13 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 13 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 13 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 89 13 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 88 13 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 88 13 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 13 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 13 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 87 13 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 86 13 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 86 13 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 85 13 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 85 13 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 13 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 13 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 84 13 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 83 13 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 13 83 13 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 13 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 13 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 13 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 81 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 81 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 13 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 13 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 13 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 79 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 79 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 13 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 13 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 13 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 77 13 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 77 13 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 76 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 76 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 13 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 13 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 13 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 74 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 74 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 13 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 13 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 13 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 72 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 72 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 13 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 13 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 13 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 70 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 70 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 13 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 13 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 13 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 68 13 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 22 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 22 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 21 13 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 21 13 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 13 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 13 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 13 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 19 13 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 19 13 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 18 13 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 18 13 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 93 12 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 92 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 92 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 91 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 91 12 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 91 12 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 90 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 90 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 89 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 89 12 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 89 12 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 88 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 88 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 87 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 87 12 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 87 12 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 86 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 86 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 85 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 85 12 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 84 12 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 84 12 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 84 12 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 83 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 83 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 12 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 12 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 81 12 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 81 12 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 12 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 12 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 12 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 79 12 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 79 12 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 12 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 12 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 12 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 77 12 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 77 12 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 76 12 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 76 12 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 12 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 12 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 12 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 74 12 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 74 12 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 12 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 12 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 12 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 72 12 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 72 12 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 12 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 12 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 12 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 70 12 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 70 12 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 12 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 12 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 12 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 68 12 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 22 12 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 22 12 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 21 12 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 21 12 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 12 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 12 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 12 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 19 12 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 19 12 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 93 12 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 92 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 92 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 91 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 91 12 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 91 12 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 90 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 90 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 89 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 89 12 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 89 12 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 88 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 88 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 87 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 87 12 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 87 12 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 86 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 86 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 85 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 85 12 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 84 12 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 84 12 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 84 12 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 83 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 83 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 12 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 82 12 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 81 12 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 81 12 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 12 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 12 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 80 12 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 79 12 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 79 12 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 12 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 12 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 78 12 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 77 12 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 77 12 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 76 12 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 76 12 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 12 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 12 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 75 12 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 74 12 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 74 12 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 12 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 12 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 73 12 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 72 12 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 72 12 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 12 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 12 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 71 12 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 70 12 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 70 12 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 12 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 12 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 69 12 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 68 12 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 22 12 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 22 12 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 21 12 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 21 12 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 12 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 12 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 20 12 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 19 12 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 19 12 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 12 18 12 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 93 12 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 92 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 92 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 12 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 12 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 12 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 90 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 90 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 12 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 12 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 12 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 88 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 88 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 12 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 12 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 12 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 86 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 86 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 85 12 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 85 12 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 12 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 12 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 12 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 83 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 83 12 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 82 11 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 82 11 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 82 11 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 81 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 81 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 80 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 80 11 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 80 11 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 79 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 79 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 78 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 78 11 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 78 11 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 77 11 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 77 11 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 76 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 76 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 75 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 75 11 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 75 11 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 74 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 74 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 73 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 73 11 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 73 11 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 72 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 72 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 71 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 71 11 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 71 11 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 70 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 70 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 69 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 69 11 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 69 11 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 68 11 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 22 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 22 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 21 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 21 11 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 20 11 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 20 11 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 20 11 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 19 11 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 19 11 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 93 11 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 92 11 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 92 11 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 11 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 11 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 11 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 90 11 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 90 11 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 11 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 11 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 11 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 88 11 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 88 11 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 11 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 11 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 11 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 86 11 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 86 11 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 85 11 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 85 11 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 11 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 11 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 11 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 83 11 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 83 11 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 82 11 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 82 11 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 82 11 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 81 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 81 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 80 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 80 11 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 80 11 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 79 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 79 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 78 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 78 11 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 78 11 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 77 11 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 77 11 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 76 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 76 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 75 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 75 11 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 75 11 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 74 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 74 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 73 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 73 11 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 73 11 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 72 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 72 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 71 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 71 11 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 71 11 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 70 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 70 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 69 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 69 11 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 69 11 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 68 11 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 22 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 22 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 21 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 21 11 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 20 11 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 20 11 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 20 11 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 19 11 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 19 11 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 18 11 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 93 11 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 92 11 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 92 11 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 11 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 11 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 91 11 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 90 11 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 90 11 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 11 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 11 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 89 11 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 88 11 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 88 11 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 11 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 11 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 87 11 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 86 11 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 86 11 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 85 11 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 85 11 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 11 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 11 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 84 11 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 83 11 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 11 83 11 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 11 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 11 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 11 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 81 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 81 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 11 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 11 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 11 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 79 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 79 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 11 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 11 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 11 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 77 11 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 77 11 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 76 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 76 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 11 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 11 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 11 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 74 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 74 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 11 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 11 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 11 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 72 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 72 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 11 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 11 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 11 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 70 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 70 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 11 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 11 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 11 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 68 11 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 22 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 22 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 21 11 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 21 11 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 11 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 11 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 11 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 19 11 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 19 11 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 18 11 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 18 11 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 93 10 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 92 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 92 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 91 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 91 10 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 91 10 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 90 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 90 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 89 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 89 10 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 89 10 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 88 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 88 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 87 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 87 10 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 87 10 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 86 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 86 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 85 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 85 10 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 84 10 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 84 10 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 84 10 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 83 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 83 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 10 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 10 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 81 10 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 81 10 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 10 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 10 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 10 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 79 10 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 79 10 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 10 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 10 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 10 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 77 10 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 77 10 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 76 10 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 76 10 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 10 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 10 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 10 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 74 10 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 74 10 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 10 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 10 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 10 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 72 10 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 72 10 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 10 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 10 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 10 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 70 10 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 70 10 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 10 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 10 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 10 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 68 10 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 22 10 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 22 10 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 21 10 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 21 10 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 10 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 10 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 10 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 19 10 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 19 10 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 93 10 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 92 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 92 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 91 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 91 10 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 91 10 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 90 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 90 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 89 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 89 10 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 89 10 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 88 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 88 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 87 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 87 10 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 87 10 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 86 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 86 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 85 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 85 10 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 84 10 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 84 10 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 84 10 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 83 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 83 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 10 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 82 10 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 81 10 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 81 10 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 10 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 10 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 80 10 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 79 10 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 79 10 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 10 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 10 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 78 10 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 77 10 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 77 10 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 76 10 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 76 10 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 10 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 10 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 75 10 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 74 10 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 74 10 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 10 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 10 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 73 10 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 72 10 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 72 10 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 10 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 10 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 71 10 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 70 10 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 70 10 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 10 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 10 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 69 10 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 68 10 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 22 10 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 22 10 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 21 10 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 21 10 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 10 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 10 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 20 10 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 19 10 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 19 10 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 10 18 10 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 93 10 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 92 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 92 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 10 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 10 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 10 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 90 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 90 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 10 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 10 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 10 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 88 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 88 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 10 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 10 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 10 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 86 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 86 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 85 10 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 85 10 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 10 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 10 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 10 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 83 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 83 10 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 82 9 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 82 9 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 82 9 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 81 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 81 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 80 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 80 9 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 80 9 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 79 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 79 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 78 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 78 9 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 78 9 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 77 9 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 77 9 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 76 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 76 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 75 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 75 9 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 75 9 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 74 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 74 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 73 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 73 9 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 73 9 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 72 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 72 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 71 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 71 9 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 71 9 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 70 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 70 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 69 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 69 9 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 69 9 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 68 9 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 22 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 22 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 21 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 21 9 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 20 9 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 20 9 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 20 9 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 19 9 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 19 9 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 93 9 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 92 9 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 92 9 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 9 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 9 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 9 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 90 9 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 90 9 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 9 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 9 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 9 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 88 9 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 88 9 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 9 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 9 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 9 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 86 9 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 86 9 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 85 9 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 85 9 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 9 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 9 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 9 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 83 9 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 83 9 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 82 9 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 82 9 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 82 9 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 81 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 81 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 80 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 80 9 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 80 9 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 79 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 79 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 78 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 78 9 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 78 9 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 77 9 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 77 9 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 76 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 76 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 75 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 75 9 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 75 9 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 74 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 74 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 73 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 73 9 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 73 9 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 72 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 72 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 71 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 71 9 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 71 9 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 70 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 70 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 69 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 69 9 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 69 9 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 68 9 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 22 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 22 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 21 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 21 9 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 20 9 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 20 9 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 20 9 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 19 9 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 19 9 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 18 9 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 93 9 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 92 9 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 92 9 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 9 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 9 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 91 9 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 90 9 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 90 9 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 9 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 9 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 89 9 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 88 9 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 88 9 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 9 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 9 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 87 9 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 86 9 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 86 9 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 85 9 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 85 9 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 9 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 9 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 84 9 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 83 9 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 9 83 9 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 9 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 9 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 9 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 81 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 81 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 9 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 9 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 9 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 79 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 79 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 9 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 9 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 9 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 77 9 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 77 9 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 76 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 76 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 9 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 9 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 9 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 74 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 74 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 9 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 9 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 9 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 72 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 72 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 9 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 9 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 9 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 70 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 70 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 9 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 9 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 9 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 68 9 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 22 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 22 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 21 9 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 21 9 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 9 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 9 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 9 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 19 9 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 19 9 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 18 9 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 18 9 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 93 8 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 92 8 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 92 8 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 91 8 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 91 8 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 91 8 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 90 8 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 90 8 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 89 8 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 89 8 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 89 8 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 88 8 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 88 8 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 87 8 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 87 8 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 87 8 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 86 8 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 86 8 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 85 8 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 85 8 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 84 8 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 84 8 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 84 8 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 83 8 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 83 8 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 8 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 8 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 8 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 81 8 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 81 8 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 8 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 8 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 8 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 79 8 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 79 8 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 8 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 8 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 8 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 77 8 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 77 8 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 76 8 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 76 8 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 8 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 8 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 8 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 74 8 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 74 8 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 8 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 8 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 8 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 72 8 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 72 8 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 8 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 8 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 8 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 70 8 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 70 8 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 8 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 8 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 8 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 68 8 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 22 8 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 22 8 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 21 8 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 21 8 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 8 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 8 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 8 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 19 8 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 19 8 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 93 8 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 92 8 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 92 8 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 91 8 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 91 8 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 91 8 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 90 8 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 90 8 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 89 8 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 89 8 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 89 8 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 88 8 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 88 8 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 87 8 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 87 8 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 87 8 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 86 8 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 86 8 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 85 8 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 85 8 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 84 8 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 84 8 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 84 8 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 83 8 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 83 8 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 8 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 8 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 82 8 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 81 8 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 81 8 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 8 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 8 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 80 8 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 79 8 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 79 8 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 8 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 8 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 78 8 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 77 8 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 77 8 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 76 8 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 76 8 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 8 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 8 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 75 8 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 74 8 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 74 8 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 8 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 8 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 73 8 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 72 8 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 72 8 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 8 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 8 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 71 8 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 70 8 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 70 8 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 8 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 8 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 69 8 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 68 8 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 22 8 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 22 8 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 21 8 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 21 8 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 8 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 8 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 20 8 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 19 8 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 19 8 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 8 18 8 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 93 7 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 92 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 92 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 91 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 91 7 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 91 7 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 90 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 90 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 89 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 89 7 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 89 7 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 88 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 88 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 87 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 87 7 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 87 7 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 86 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 86 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 85 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 85 7 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 84 7 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 84 7 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 84 7 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 83 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 83 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 82 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 82 7 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 82 7 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 81 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 81 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 80 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 80 7 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 80 7 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 79 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 79 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 78 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 78 7 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 78 7 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 77 7 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 77 7 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 76 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 76 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 75 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 75 7 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 75 7 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 74 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 74 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 73 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 73 7 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 73 7 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 72 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 72 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 71 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 71 7 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 71 7 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 70 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 70 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 69 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 69 7 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 69 7 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 68 7 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 22 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 22 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 21 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 21 7 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 20 7 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 20 7 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 20 7 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 19 7 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 19 7 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 93 7 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 92 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 92 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 91 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 91 7 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 91 7 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 90 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 90 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 89 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 89 7 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 89 7 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 88 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 88 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 87 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 87 7 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 87 7 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 86 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 86 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 85 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 85 7 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 84 7 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 84 7 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 84 7 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 83 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 83 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 82 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 82 7 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 82 7 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 81 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 81 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 80 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 80 7 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 80 7 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 79 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 79 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 78 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 78 7 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 78 7 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 77 7 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 77 7 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 76 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 76 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 75 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 75 7 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 75 7 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 74 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 74 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 73 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 73 7 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 73 7 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 72 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 72 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 71 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 71 7 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 71 7 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 70 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 70 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 69 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 69 7 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 69 7 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 68 7 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 22 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 22 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 21 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 21 7 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 20 7 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 20 7 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 20 7 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 19 7 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 19 7 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 7 18 7 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 93 7 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 92 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 92 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 7 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 7 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 7 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 90 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 90 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 7 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 7 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 7 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 88 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 88 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 7 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 7 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 7 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 86 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 86 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 85 7 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 85 7 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 7 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 7 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 7 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 83 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 83 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 7 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 7 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 7 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 81 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 81 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 7 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 7 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 7 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 79 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 79 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 7 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 7 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 7 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 77 7 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 77 7 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 76 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 76 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 7 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 7 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 7 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 74 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 74 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 7 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 7 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 7 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 72 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 72 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 7 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 7 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 7 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 70 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 70 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 7 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 7 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 7 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 68 7 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 22 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 22 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 21 7 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 21 7 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 7 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 7 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 7 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 19 7 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 19 7 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 18 7 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 18 7 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 93 6 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 92 6 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 92 6 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 6 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 6 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 6 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 90 6 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 90 6 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 6 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 6 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 6 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 88 6 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 88 6 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 6 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 6 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 6 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 86 6 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 86 6 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 85 6 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 85 6 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 6 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 6 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 6 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 83 6 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 83 6 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 6 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 6 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 6 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 81 6 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 81 6 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 6 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 6 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 6 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 79 6 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 79 6 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 6 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 6 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 6 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 77 6 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 77 6 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 76 6 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 76 6 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 6 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 6 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 6 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 74 6 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 74 6 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 6 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 6 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 6 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 72 6 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 72 6 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 6 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 6 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 6 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 70 6 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 70 6 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 6 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 6 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 6 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 68 6 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 22 6 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 22 6 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 21 6 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 21 6 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 6 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 6 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 6 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 19 6 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 19 6 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 93 6 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 92 6 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 92 6 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 6 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 6 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 91 6 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 90 6 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 90 6 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 6 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 6 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 89 6 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 88 6 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 88 6 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 6 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 6 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 87 6 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 86 6 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 86 6 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 85 6 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 85 6 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 6 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 6 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 84 6 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 83 6 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 83 6 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 6 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 6 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 82 6 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 81 6 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 81 6 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 6 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 6 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 80 6 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 79 6 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 79 6 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 6 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 6 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 78 6 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 77 6 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 77 6 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 76 6 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 76 6 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 6 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 6 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 75 6 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 74 6 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 74 6 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 6 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 6 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 73 6 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 72 6 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 72 6 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 6 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 6 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 71 6 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 70 6 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 70 6 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 6 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 6 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 69 6 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 68 6 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 22 6 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 22 6 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 21 6 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 21 6 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 6 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 6 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 20 6 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 19 6 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 19 6 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 6 18 6 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 93 5 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 92 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 92 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 91 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 91 5 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 91 5 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 90 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 90 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 89 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 89 5 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 89 5 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 88 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 88 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 87 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 87 5 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 87 5 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 86 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 86 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 85 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 85 5 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 84 5 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 84 5 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 84 5 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 83 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 83 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 82 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 82 5 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 82 5 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 81 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 81 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 80 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 80 5 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 80 5 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 79 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 79 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 78 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 78 5 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 78 5 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 77 5 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 77 5 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 76 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 76 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 75 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 75 5 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 75 5 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 74 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 74 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 73 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 73 5 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 73 5 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 72 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 72 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 71 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 71 5 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 71 5 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 70 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 70 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 69 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 69 5 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 69 5 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 68 5 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 22 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 22 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 21 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 21 5 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 20 5 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 20 5 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 20 5 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 19 5 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 19 5 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 82 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 82 5 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 82 5 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 81 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 81 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 80 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 80 5 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 80 5 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 79 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 79 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 78 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 78 5 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 78 5 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 77 5 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 77 5 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 76 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 76 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 75 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 75 5 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 75 5 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 74 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 74 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 73 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 73 5 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 73 5 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 72 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 72 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 71 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 71 5 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 71 5 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 70 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 70 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 69 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 69 5 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 69 5 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 68 5 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 93 5 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 92 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 92 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 91 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 91 5 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 91 5 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 90 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 90 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 89 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 89 5 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 89 5 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 88 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 88 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 87 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 87 5 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 87 5 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 86 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 86 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 85 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 85 5 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 84 5 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 84 5 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 84 5 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 83 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 83 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 22 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 22 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 21 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 21 5 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 20 5 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 20 5 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 20 5 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 19 5 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 19 5 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 5 18 5 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 5 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 5 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 81 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 81 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 5 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 5 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 5 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 79 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 79 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 5 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 5 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 5 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 77 5 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 77 5 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 76 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 76 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 5 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 5 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 5 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 74 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 74 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 5 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 5 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 5 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 72 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 72 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 5 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 5 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 5 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 70 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 70 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 5 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 5 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 5 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 68 5 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 93 5 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 92 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 92 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 5 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 5 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 5 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 90 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 90 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 5 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 5 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 5 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 88 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 88 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 5 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 5 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 5 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 86 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 86 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 85 5 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 85 5 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 5 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 5 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 5 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 83 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 83 5 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 22 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 22 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 21 5 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 21 5 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 5 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 5 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 5 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 19 5 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 19 5 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 18 5 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 18 5 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 4 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 4 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 4 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 81 4 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 81 4 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 4 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 4 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 4 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 79 4 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 79 4 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 4 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 4 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 4 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 77 4 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 77 4 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 76 4 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 76 4 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 4 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 4 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 4 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 74 4 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 74 4 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 4 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 4 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 4 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 72 4 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 72 4 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 4 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 4 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 4 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 70 4 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 70 4 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 4 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 4 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 4 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 68 4 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 93 4 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 92 4 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 92 4 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 4 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 4 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 4 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 90 4 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 90 4 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 4 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 4 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 4 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 88 4 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 88 4 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 4 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 4 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 4 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 86 4 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 86 4 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 85 4 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 85 4 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 4 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 4 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 4 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 83 4 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 83 4 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 22 4 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 22 4 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 21 4 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 21 4 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 4 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 4 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 4 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 19 4 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 19 4 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 4 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 4 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 82 4 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 81 4 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 81 4 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 4 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 4 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 80 4 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 79 4 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 79 4 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 4 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 4 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 78 4 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 77 4 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 77 4 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 76 4 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 76 4 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 4 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 4 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 75 4 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 74 4 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 74 4 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 4 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 4 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 73 4 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 72 4 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 72 4 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 4 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 4 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 71 4 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 70 4 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 70 4 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 4 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 4 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 69 4 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 68 4 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 93 4 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 92 4 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 92 4 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 4 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 4 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 91 4 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 90 4 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 90 4 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 4 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 4 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 89 4 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 88 4 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 88 4 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 4 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 4 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 87 4 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 86 4 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 86 4 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 85 4 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 85 4 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 4 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 4 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 84 4 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 83 4 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 83 4 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 22 4 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 22 4 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 21 4 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 21 4 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 4 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 4 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 20 4 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 19 4 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 19 4 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 4 18 4 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 82 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 82 3 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 82 3 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 81 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 81 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 80 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 80 3 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 80 3 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 79 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 79 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 78 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 78 3 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 78 3 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 77 3 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 77 3 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 76 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 76 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 75 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 75 3 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 75 3 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 74 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 74 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 73 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 73 3 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 73 3 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 72 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 72 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 71 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 71 3 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 71 3 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 70 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 70 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 69 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 69 3 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 69 3 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 68 3 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 93 3 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 92 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 92 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 91 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 91 3 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 91 3 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 90 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 90 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 89 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 89 3 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 89 3 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 88 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 88 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 87 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 87 3 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 87 3 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 86 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 86 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 85 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 85 3 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 84 3 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 84 3 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 84 3 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 83 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 83 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 22 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 22 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 21 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 21 3 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 20 3 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 20 3 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 20 3 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 19 3 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 19 3 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 82 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 82 3 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 82 3 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 81 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 81 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 80 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 80 3 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 80 3 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 79 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 79 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 78 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 78 3 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 78 3 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 77 3 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 77 3 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 76 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 76 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 75 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 75 3 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 75 3 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 74 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 74 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 73 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 73 3 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 73 3 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 72 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 72 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 71 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 71 3 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 71 3 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 70 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 70 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 69 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 69 3 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 69 3 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 68 3 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 93 3 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 92 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 92 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 91 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 91 3 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 91 3 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 90 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 90 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 89 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 89 3 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 89 3 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 88 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 88 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 87 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 87 3 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 87 3 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 86 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 86 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 85 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 85 3 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 84 3 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 84 3 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 84 3 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 83 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 83 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 22 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 22 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 21 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 21 3 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 20 3 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 20 3 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 20 3 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 19 3 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 19 3 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 3 18 3 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 3 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 3 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 81 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 81 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 3 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 3 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 3 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 79 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 79 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 3 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 3 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 3 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 77 3 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 77 3 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 76 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 76 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 3 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 3 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 3 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 74 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 74 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 3 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 3 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 3 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 72 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 72 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 3 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 3 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 3 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 70 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 70 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 3 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 3 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 3 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 68 3 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 93 3 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 92 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 92 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 3 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 3 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 3 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 90 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 90 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 3 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 3 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 3 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 88 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 88 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 3 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 3 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 3 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 86 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 86 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 85 3 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 85 3 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 3 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 3 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 3 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 83 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 83 3 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 22 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 22 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 21 3 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 21 3 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 3 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 3 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 3 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 19 3 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 19 3 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 18 3 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 18 3 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 2 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 2 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 2 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 81 2 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 81 2 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 2 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 2 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 2 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 79 2 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 79 2 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 2 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 2 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 2 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 77 2 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 77 2 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 76 2 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 76 2 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 2 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 2 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 2 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 74 2 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 74 2 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 2 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 2 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 2 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 72 2 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 72 2 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 2 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 2 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 2 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 70 2 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 70 2 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 2 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 2 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 2 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 68 2 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 93 2 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 92 2 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 92 2 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 2 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 2 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 2 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 90 2 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 90 2 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 2 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 2 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 2 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 88 2 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 88 2 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 2 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 2 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 2 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 86 2 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 86 2 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 85 2 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 85 2 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 2 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 2 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 2 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 83 2 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 83 2 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 22 2 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 22 2 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 21 2 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 21 2 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 2 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 2 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 2 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 19 2 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 19 2 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 2 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 2 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 82 2 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 81 2 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 81 2 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 2 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 2 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 80 2 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 79 2 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 79 2 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 2 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 2 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 78 2 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 77 2 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 77 2 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 76 2 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 76 2 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 2 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 2 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 75 2 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 74 2 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 74 2 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 2 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 2 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 73 2 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 72 2 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 72 2 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 2 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 2 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 71 2 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 70 2 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 70 2 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 2 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 2 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 69 2 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 68 2 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 93 2 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 92 2 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 92 2 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 2 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 2 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 91 2 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 90 2 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 90 2 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 2 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 2 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 89 2 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 88 2 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 88 2 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 2 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 2 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 87 2 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 86 2 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 86 2 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 85 2 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 85 2 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 2 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 2 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 84 2 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 83 2 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 83 2 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 22 2 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 22 2 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 21 2 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 21 2 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 2 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 2 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 20 2 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 19 2 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 19 2 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 2 18 2 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 82 1 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 82 1 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 82 1 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 81 1 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 81 1 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 80 1 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 80 1 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 80 1 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 79 1 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 79 1 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 78 1 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 78 1 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 78 1 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 77 1 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 77 1 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 76 1 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 76 1 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 75 1 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 75 1 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 75 1 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 74 1 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 74 1 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 73 1 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 73 1 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 73 1 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 72 1 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 72 1 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 71 1 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 71 1 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 71 1 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 70 1 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 70 1 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 69 1 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 69 1 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 69 1 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 68 1 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 93 1 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 92 1 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 92 1 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 91 1 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 91 1 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 91 1 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 90 1 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 90 1 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 89 1 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 89 1 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 89 1 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 88 1 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 88 1 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 87 1 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 87 1 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 87 1 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 86 1 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 86 1 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 85 1 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 85 1 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 84 1 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 84 1 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 84 1 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 83 1 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 83 1 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 22 1 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 22 1 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 21 1 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 21 1 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 20 1 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 20 1 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 20 1 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 19 1 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 19 1 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 82 1 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 82 1 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 82 1 82 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 81 1 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 81 1 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 80 1 81 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 80 1 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 80 1 80 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 79 1 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 79 1 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 78 1 79 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 78 1 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 78 1 78 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 77 1 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 77 1 77 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 76 1 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 76 1 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 75 1 76 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 75 1 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 75 1 75 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 74 1 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 74 1 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 73 1 74 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 73 1 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 73 1 73 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 72 1 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 72 1 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 71 1 72 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 71 1 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 71 1 71 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 70 1 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 70 1 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 69 1 70 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 69 1 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 69 1 69 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 68 1 68 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 93 1 93 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 92 1 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 92 1 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 91 1 92 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 91 1 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 91 1 91 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 90 1 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 90 1 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 89 1 90 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 89 1 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 89 1 89 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 88 1 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 88 1 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 87 1 88 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 87 1 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 87 1 87 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 86 1 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 86 1 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 85 1 86 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 85 1 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 84 1 85 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 84 1 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 84 1 84 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 83 1 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 83 1 83 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 22 1 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 22 1 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 21 1 22 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 21 1 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 20 1 21 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 20 1 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 20 1 20 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 19 1 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 19 1 19 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDIO
port 6 nsew power bidirectional
rlabel nfet_brown s 1 18 1 18 6 VDDIO
port 6 nsew power bidirectional
rlabel 
 s 1 62 25 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel 
 s 51 62 75 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 62 24 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 51 62 75 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 66 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 66 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 75 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 75 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 64 75 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 64 75 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 75 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 75 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 75 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 62 75 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 66 74 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 66 74 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 74 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 74 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 74 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 64 74 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 64 74 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 74 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 74 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 74 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 62 74 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 66 74 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 66 74 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 74 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 74 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 65 74 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 64 74 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 64 74 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 74 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 74 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 63 74 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 74 62 74 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 66 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 66 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 65 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 65 73 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 65 73 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 64 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 64 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 63 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 63 73 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 63 73 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 62 73 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 66 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 66 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 65 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 65 73 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 65 73 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 64 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 64 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 63 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 63 73 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 63 73 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 73 62 73 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 66 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 66 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 73 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 73 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 73 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 64 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 64 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 73 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 73 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 73 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 62 73 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 66 72 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 66 72 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 72 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 72 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 72 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 64 72 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 64 72 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 72 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 72 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 72 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 62 72 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 66 72 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 66 72 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 72 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 72 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 65 72 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 64 72 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 64 72 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 72 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 72 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 63 72 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 72 62 72 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 66 71 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 66 71 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 65 71 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 65 71 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 65 71 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 64 71 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 64 71 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 63 71 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 63 71 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 63 71 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 62 71 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 66 71 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 66 71 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 65 71 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 65 71 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 65 71 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 64 71 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 64 71 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 63 71 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 63 71 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 63 71 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 71 62 71 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 66 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 66 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 65 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 65 70 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 65 70 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 64 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 64 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 63 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 63 70 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 63 70 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 62 70 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 66 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 66 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 65 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 65 70 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 65 70 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 64 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 64 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 63 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 63 70 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 63 70 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 70 62 70 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 66 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 66 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 70 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 70 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 70 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 64 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 64 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 70 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 70 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 70 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 62 70 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 66 69 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 66 69 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 69 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 69 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 69 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 64 69 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 64 69 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 69 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 69 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 69 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 62 69 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 66 69 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 66 69 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 69 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 69 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 65 69 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 64 69 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 64 69 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 69 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 69 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 63 69 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 69 62 69 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 66 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 66 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 65 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 65 68 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 65 68 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 64 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 64 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 63 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 63 68 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 63 68 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 62 68 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 66 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 66 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 65 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 65 68 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 65 68 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 64 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 64 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 63 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 63 68 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 63 68 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 68 62 68 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 66 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 66 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 68 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 68 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 68 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 64 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 64 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 68 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 68 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 68 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 62 68 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 66 67 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 66 67 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 67 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 67 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 67 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 64 67 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 64 67 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 67 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 67 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 67 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 62 67 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 66 67 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 66 67 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 67 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 67 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 65 67 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 64 67 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 64 67 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 67 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 67 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 63 67 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 67 62 67 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 66 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 66 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 65 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 65 66 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 65 66 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 64 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 64 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 63 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 63 66 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 63 66 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 62 66 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 66 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 66 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 65 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 65 66 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 65 66 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 64 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 64 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 63 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 63 66 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 63 66 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 66 62 66 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 66 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 66 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 66 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 66 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 66 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 64 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 64 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 66 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 66 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 66 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 62 66 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 66 65 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 66 65 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 65 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 65 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 65 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 64 65 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 64 65 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 65 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 65 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 65 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 62 65 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 66 65 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 66 65 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 65 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 65 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 65 65 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 64 65 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 64 65 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 65 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 65 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 63 65 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 65 62 65 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 66 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 66 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 65 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 65 64 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 65 64 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 64 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 64 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 63 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 63 64 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 63 64 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 62 64 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 66 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 66 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 65 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 65 64 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 65 64 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 64 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 64 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 63 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 63 64 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 63 64 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 64 62 64 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 66 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 66 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 64 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 64 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 64 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 64 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 64 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 64 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 64 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 64 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 62 64 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 66 63 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 66 63 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 63 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 63 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 63 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 64 63 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 64 63 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 63 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 63 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 63 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 62 63 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 66 63 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 66 63 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 63 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 63 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 65 63 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 64 63 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 64 63 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 63 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 63 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 63 63 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 63 62 63 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 66 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 66 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 65 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 65 62 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 65 62 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 64 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 64 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 63 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 63 62 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 63 62 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 62 62 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 66 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 66 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 65 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 65 62 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 65 62 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 64 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 64 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 63 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 63 62 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 63 62 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 62 62 62 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 66 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 66 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 62 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 62 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 62 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 64 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 64 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 62 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 62 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 62 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 62 62 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 66 61 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 66 61 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 61 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 61 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 61 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 64 61 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 64 61 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 61 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 61 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 61 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 62 61 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 66 61 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 66 61 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 61 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 61 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 65 61 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 64 61 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 64 61 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 61 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 61 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 63 61 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 61 62 61 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 66 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 66 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 65 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 65 60 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 65 60 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 64 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 64 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 63 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 63 60 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 63 60 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 62 60 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 66 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 66 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 65 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 65 60 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 65 60 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 64 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 64 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 63 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 63 60 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 63 60 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 60 62 60 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 66 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 66 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 60 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 60 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 60 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 64 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 64 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 60 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 60 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 60 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 62 60 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 66 59 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 66 59 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 59 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 59 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 59 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 64 59 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 64 59 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 59 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 59 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 59 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 62 59 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 66 59 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 66 59 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 59 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 59 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 65 59 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 64 59 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 64 59 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 59 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 59 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 63 59 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 59 62 59 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 66 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 66 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 65 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 65 58 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 65 58 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 64 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 64 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 63 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 63 58 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 63 58 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 62 58 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 66 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 66 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 65 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 65 58 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 65 58 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 64 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 64 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 63 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 63 58 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 63 58 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 58 62 58 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 66 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 66 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 58 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 58 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 58 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 64 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 64 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 58 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 58 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 58 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 62 58 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 66 57 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 66 57 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 57 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 57 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 57 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 64 57 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 64 57 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 57 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 57 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 57 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 62 57 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 66 57 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 66 57 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 57 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 57 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 65 57 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 64 57 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 64 57 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 57 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 57 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 63 57 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 57 62 57 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 66 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 66 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 65 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 65 56 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 65 56 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 64 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 64 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 63 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 63 56 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 63 56 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 62 56 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 66 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 66 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 65 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 65 56 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 65 56 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 64 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 64 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 63 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 63 56 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 63 56 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 56 62 56 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 66 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 66 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 65 56 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 65 56 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 65 56 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 64 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 64 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 63 56 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 63 56 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 63 56 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 62 56 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 66 55 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 66 55 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 65 55 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 65 55 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 65 55 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 64 55 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 64 55 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 63 55 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 63 55 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 63 55 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 55 62 55 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 66 55 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 66 55 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 55 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 55 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 55 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 64 55 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 64 55 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 55 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 55 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 55 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 62 55 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 66 54 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 66 54 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 54 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 54 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 54 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 64 54 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 64 54 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 54 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 54 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 54 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 62 54 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 66 54 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 66 54 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 54 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 54 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 65 54 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 64 54 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 64 54 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 54 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 54 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 63 54 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 54 62 54 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 66 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 66 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 65 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 65 53 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 65 53 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 64 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 64 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 63 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 63 53 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 63 53 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 62 53 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 66 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 66 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 65 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 65 53 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 65 53 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 64 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 64 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 63 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 63 53 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 63 53 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 53 62 53 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 66 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 66 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 53 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 53 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 53 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 64 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 64 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 53 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 53 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 53 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 62 53 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 66 52 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 66 52 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 52 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 52 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 52 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 64 52 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 64 52 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 52 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 52 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 52 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 62 52 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 66 52 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 66 52 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 52 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 52 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 65 52 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 64 52 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 64 52 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 52 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 52 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 63 52 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 52 62 52 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 66 51 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 66 51 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 65 51 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 65 51 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 65 51 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 64 51 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 64 51 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 63 51 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 63 51 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 63 51 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 62 51 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 66 51 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 66 51 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 65 51 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 65 51 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 65 51 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 64 51 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 64 51 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 63 51 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 63 51 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 63 51 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 51 62 51 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 66 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 66 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 65 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 65 24 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 65 24 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 64 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 64 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 63 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 63 24 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 63 24 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 62 24 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 66 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 66 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 65 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 65 24 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 65 24 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 64 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 64 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 63 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 63 24 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 63 24 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 24 62 24 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 66 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 66 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 24 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 24 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 24 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 64 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 64 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 24 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 24 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 24 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 62 24 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 66 23 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 66 23 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 23 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 23 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 23 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 64 23 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 64 23 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 23 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 23 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 23 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 62 23 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 66 23 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 66 23 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 23 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 23 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 65 23 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 64 23 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 64 23 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 23 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 23 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 63 23 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 23 62 23 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 66 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 66 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 65 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 65 22 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 65 22 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 64 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 64 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 63 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 63 22 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 63 22 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 62 22 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 66 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 66 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 65 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 65 22 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 65 22 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 64 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 64 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 63 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 63 22 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 63 22 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 22 62 22 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 66 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 66 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 22 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 22 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 22 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 64 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 64 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 22 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 22 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 22 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 62 22 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 66 21 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 66 21 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 21 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 21 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 21 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 64 21 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 64 21 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 21 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 21 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 21 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 62 21 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 66 21 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 66 21 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 21 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 21 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 65 21 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 64 21 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 64 21 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 21 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 21 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 63 21 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 21 62 21 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 66 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 66 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 65 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 65 20 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 65 20 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 64 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 64 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 63 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 63 20 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 63 20 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 62 20 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 66 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 66 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 65 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 65 20 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 65 20 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 64 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 64 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 63 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 63 20 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 63 20 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 20 62 20 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 66 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 66 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 20 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 20 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 20 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 64 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 64 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 20 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 20 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 20 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 62 20 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 66 19 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 66 19 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 19 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 19 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 19 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 64 19 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 64 19 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 19 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 19 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 19 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 62 19 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 66 19 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 66 19 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 19 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 19 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 65 19 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 64 19 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 64 19 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 19 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 19 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 63 19 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 19 62 19 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 66 18 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 66 18 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 65 18 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 65 18 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 65 18 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 64 18 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 64 18 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 63 18 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 63 18 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 63 18 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 62 18 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 66 18 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 66 18 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 65 18 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 65 18 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 65 18 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 64 18 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 64 18 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 63 18 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 63 18 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 63 18 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 18 62 18 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 66 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 66 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 65 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 65 17 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 65 17 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 64 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 64 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 63 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 63 17 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 63 17 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 62 17 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 66 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 66 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 65 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 65 17 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 65 17 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 64 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 64 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 63 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 63 17 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 63 17 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 17 62 17 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 66 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 66 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 17 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 17 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 17 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 64 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 64 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 17 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 17 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 17 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 62 17 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 66 16 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 66 16 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 16 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 16 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 16 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 64 16 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 64 16 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 16 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 16 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 16 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 62 16 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 66 16 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 66 16 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 16 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 16 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 65 16 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 64 16 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 64 16 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 16 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 16 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 63 16 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 16 62 16 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 66 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 66 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 65 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 65 15 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 65 15 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 64 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 64 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 63 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 63 15 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 63 15 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 62 15 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 66 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 66 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 65 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 65 15 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 65 15 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 64 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 64 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 63 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 63 15 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 63 15 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 15 62 15 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 66 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 66 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 15 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 15 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 15 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 64 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 64 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 15 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 15 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 15 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 62 15 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 66 14 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 66 14 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 14 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 14 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 14 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 64 14 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 64 14 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 14 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 14 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 14 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 62 14 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 66 14 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 66 14 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 14 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 14 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 65 14 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 64 14 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 64 14 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 14 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 14 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 63 14 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 14 62 14 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 66 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 66 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 65 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 65 13 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 65 13 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 64 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 64 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 63 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 63 13 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 63 13 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 62 13 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 66 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 66 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 65 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 65 13 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 65 13 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 64 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 64 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 63 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 63 13 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 63 13 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 13 62 13 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 66 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 66 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 13 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 13 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 13 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 64 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 64 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 13 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 13 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 13 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 62 13 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 66 12 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 66 12 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 12 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 12 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 12 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 64 12 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 64 12 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 12 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 12 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 12 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 62 12 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 66 12 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 66 12 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 12 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 12 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 65 12 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 64 12 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 64 12 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 12 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 12 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 63 12 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 12 62 12 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 66 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 66 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 65 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 65 11 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 65 11 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 64 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 64 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 63 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 63 11 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 63 11 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 62 11 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 66 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 66 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 65 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 65 11 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 65 11 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 64 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 64 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 63 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 63 11 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 63 11 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 11 62 11 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 66 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 66 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 11 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 11 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 11 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 64 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 64 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 11 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 11 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 11 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 62 11 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 66 10 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 66 10 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 10 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 10 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 10 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 64 10 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 64 10 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 10 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 10 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 10 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 62 10 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 66 10 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 66 10 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 10 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 10 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 65 10 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 64 10 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 64 10 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 10 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 10 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 63 10 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 10 62 10 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 66 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 66 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 65 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 65 9 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 65 9 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 64 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 64 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 63 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 63 9 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 63 9 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 62 9 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 66 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 66 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 65 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 65 9 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 65 9 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 64 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 64 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 63 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 63 9 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 63 9 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 9 62 9 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 66 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 66 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 9 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 9 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 9 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 64 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 64 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 9 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 9 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 9 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 62 9 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 66 8 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 66 8 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 8 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 8 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 8 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 64 8 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 64 8 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 8 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 8 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 8 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 62 8 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 66 8 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 66 8 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 8 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 8 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 65 8 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 64 8 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 64 8 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 8 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 8 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 63 8 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 8 62 8 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 66 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 66 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 65 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 65 7 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 65 7 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 64 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 64 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 63 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 63 7 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 63 7 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 62 7 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 66 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 66 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 65 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 65 7 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 65 7 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 64 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 64 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 63 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 63 7 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 63 7 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 7 62 7 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 66 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 66 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 7 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 7 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 7 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 64 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 64 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 7 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 7 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 7 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 62 7 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 66 6 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 66 6 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 6 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 6 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 6 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 64 6 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 64 6 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 6 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 6 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 6 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 62 6 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 66 6 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 66 6 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 6 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 6 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 65 6 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 64 6 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 64 6 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 6 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 6 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 63 6 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 6 62 6 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 66 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 66 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 65 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 65 5 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 65 5 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 64 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 64 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 63 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 63 5 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 63 5 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 62 5 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 66 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 66 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 65 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 65 5 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 65 5 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 64 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 64 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 63 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 63 5 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 63 5 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 5 62 5 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 66 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 66 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 5 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 5 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 5 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 64 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 64 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 5 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 5 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 5 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 62 5 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 66 4 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 66 4 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 4 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 4 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 4 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 64 4 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 64 4 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 4 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 4 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 4 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 62 4 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 66 4 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 66 4 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 4 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 4 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 65 4 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 64 4 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 64 4 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 4 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 4 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 63 4 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 4 62 4 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 66 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 66 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 65 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 65 3 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 65 3 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 64 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 64 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 63 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 63 3 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 63 3 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 62 3 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 66 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 66 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 65 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 65 3 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 65 3 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 64 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 64 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 63 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 63 3 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 63 3 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 3 62 3 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 66 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 66 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 3 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 3 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 3 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 64 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 64 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 3 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 3 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 3 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 62 3 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 66 2 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 66 2 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 2 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 2 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 2 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 64 2 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 64 2 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 2 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 2 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 2 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 62 2 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 66 2 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 66 2 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 2 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 2 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 65 2 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 64 2 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 64 2 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 2 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 2 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 63 2 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 2 62 2 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 66 1 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 66 1 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 65 1 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 65 1 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 65 1 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 64 1 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 64 1 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 63 1 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 63 1 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 63 1 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 62 1 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 66 1 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 66 1 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 65 1 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 65 1 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 65 1 65 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 64 1 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 64 1 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 63 1 64 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 63 1 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 63 1 63 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel nfet_brown s 1 62 1 62 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 46 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 54 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 198
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
