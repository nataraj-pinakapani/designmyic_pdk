magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 11 217 277 283
rect 11 43 1052 217
rect -26 -43 1082 43
<< mvnmos >>
rect 94 107 194 257
rect 273 107 373 191
rect 415 107 515 191
rect 571 107 671 191
rect 713 107 813 191
rect 869 107 969 191
<< mvpmos >>
rect 94 443 194 743
rect 273 491 373 575
rect 415 491 515 575
rect 571 491 671 575
rect 713 491 813 575
rect 869 491 969 575
<< mvndiff >>
rect 37 249 94 257
rect 37 215 49 249
rect 83 215 94 249
rect 37 149 94 215
rect 37 115 49 149
rect 83 115 94 149
rect 37 107 94 115
rect 194 235 251 257
rect 194 201 205 235
rect 239 201 251 235
rect 194 191 251 201
rect 194 149 273 191
rect 194 115 205 149
rect 239 115 273 149
rect 194 107 273 115
rect 373 107 415 191
rect 515 166 571 191
rect 515 132 526 166
rect 560 132 571 166
rect 515 107 571 132
rect 671 107 713 191
rect 813 166 869 191
rect 813 132 824 166
rect 858 132 869 166
rect 813 107 869 132
rect 969 166 1026 191
rect 969 132 980 166
rect 1014 132 1026 166
rect 969 107 1026 132
<< mvpdiff >>
rect 37 735 94 743
rect 37 701 49 735
rect 83 701 94 735
rect 37 652 94 701
rect 37 618 49 652
rect 83 618 94 652
rect 37 568 94 618
rect 37 534 49 568
rect 83 534 94 568
rect 37 485 94 534
rect 37 451 49 485
rect 83 451 94 485
rect 37 443 94 451
rect 194 735 251 743
rect 194 701 205 735
rect 239 701 251 735
rect 194 652 251 701
rect 194 618 205 652
rect 239 618 251 652
rect 194 575 251 618
rect 194 568 273 575
rect 194 534 205 568
rect 239 534 273 568
rect 194 491 273 534
rect 373 491 415 575
rect 515 550 571 575
rect 515 516 526 550
rect 560 516 571 550
rect 515 491 571 516
rect 671 491 713 575
rect 813 550 869 575
rect 813 516 824 550
rect 858 516 869 550
rect 813 491 869 516
rect 969 550 1026 575
rect 969 516 980 550
rect 1014 516 1026 550
rect 969 491 1026 516
rect 194 485 251 491
rect 194 451 205 485
rect 239 451 251 485
rect 194 443 251 451
<< mvndiffc >>
rect 49 215 83 249
rect 49 115 83 149
rect 205 201 239 235
rect 205 115 239 149
rect 526 132 560 166
rect 824 132 858 166
rect 980 132 1014 166
<< mvpdiffc >>
rect 49 701 83 735
rect 49 618 83 652
rect 49 534 83 568
rect 49 451 83 485
rect 205 701 239 735
rect 205 618 239 652
rect 205 534 239 568
rect 526 516 560 550
rect 824 516 858 550
rect 980 516 1014 550
rect 205 451 239 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
<< poly >>
rect 94 743 194 769
rect 273 575 373 601
rect 415 575 515 601
rect 571 575 671 601
rect 713 575 813 601
rect 869 575 969 601
rect 273 443 373 491
rect 94 333 194 443
rect 94 299 140 333
rect 174 299 194 333
rect 94 257 194 299
rect 273 409 303 443
rect 337 409 373 443
rect 273 375 373 409
rect 415 469 515 491
rect 415 443 529 469
rect 415 409 475 443
rect 509 409 529 443
rect 415 393 529 409
rect 273 341 303 375
rect 337 341 373 375
rect 571 375 671 491
rect 571 351 617 375
rect 273 191 373 341
rect 423 341 617 351
rect 651 341 671 375
rect 423 321 671 341
rect 713 465 813 491
rect 713 359 819 465
rect 869 443 969 491
rect 869 409 889 443
rect 923 409 969 443
rect 869 375 969 409
rect 713 339 827 359
rect 415 217 523 321
rect 713 305 773 339
rect 807 305 827 339
rect 571 263 671 279
rect 571 229 617 263
rect 651 229 671 263
rect 415 191 515 217
rect 571 191 671 229
rect 713 271 827 305
rect 713 237 773 271
rect 807 237 827 271
rect 713 217 827 237
rect 869 341 889 375
rect 923 341 969 375
rect 713 191 813 217
rect 869 191 969 341
rect 94 81 194 107
rect 273 81 373 107
rect 415 81 515 107
rect 571 81 671 107
rect 713 81 813 107
rect 869 81 969 107
<< polycont >>
rect 140 299 174 333
rect 303 409 337 443
rect 475 409 509 443
rect 303 341 337 375
rect 617 341 651 375
rect 889 409 923 443
rect 773 305 807 339
rect 617 229 651 263
rect 773 237 807 271
rect 889 341 923 375
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 25 735 99 751
rect 25 701 49 735
rect 83 701 99 735
rect 25 652 99 701
rect 25 618 49 652
rect 83 618 99 652
rect 25 568 99 618
rect 25 534 49 568
rect 83 534 99 568
rect 25 485 99 534
rect 25 451 49 485
rect 83 451 99 485
rect 25 385 99 451
rect 135 735 251 751
rect 135 701 140 735
rect 174 701 205 735
rect 246 701 251 735
rect 135 652 251 701
rect 682 735 944 741
rect 682 701 688 735
rect 722 701 760 735
rect 794 701 832 735
rect 866 701 904 735
rect 938 701 944 735
rect 135 618 205 652
rect 239 618 251 652
rect 135 568 251 618
rect 135 534 205 568
rect 239 534 251 568
rect 135 485 251 534
rect 135 451 205 485
rect 239 451 251 485
rect 135 435 251 451
rect 287 619 646 653
rect 287 443 353 619
rect 510 550 576 583
rect 510 517 526 550
rect 287 409 303 443
rect 337 409 353 443
rect 25 249 83 385
rect 287 375 353 409
rect 124 333 190 349
rect 287 341 303 375
rect 337 341 353 375
rect 389 516 526 517
rect 560 516 576 550
rect 389 483 576 516
rect 124 299 140 333
rect 174 305 190 333
rect 389 305 423 483
rect 612 461 646 619
rect 682 550 944 701
rect 682 516 824 550
rect 858 516 944 550
rect 682 499 944 516
rect 980 550 1030 583
rect 1014 516 1030 550
rect 459 443 525 447
rect 459 409 475 443
rect 509 409 525 443
rect 612 443 935 461
rect 612 427 889 443
rect 459 391 525 409
rect 873 409 889 427
rect 923 409 935 443
rect 459 357 581 391
rect 174 299 511 305
rect 124 271 511 299
rect 25 215 49 249
rect 25 149 83 215
rect 25 115 49 149
rect 25 99 83 115
rect 119 201 205 235
rect 239 201 441 235
rect 119 149 441 201
rect 119 115 205 149
rect 239 115 441 149
rect 119 113 441 115
rect 153 79 191 113
rect 225 79 263 113
rect 297 79 335 113
rect 369 79 407 113
rect 477 183 511 271
rect 547 278 581 357
rect 617 375 737 391
rect 651 341 737 375
rect 873 375 935 409
rect 617 314 737 341
rect 773 339 823 355
rect 807 305 823 339
rect 873 341 889 375
rect 923 341 935 375
rect 873 310 935 341
rect 547 263 737 278
rect 547 229 617 263
rect 651 229 737 263
rect 547 219 737 229
rect 773 271 823 305
rect 807 255 823 271
rect 980 255 1030 516
rect 807 237 1030 255
rect 773 221 1030 237
rect 477 166 576 183
rect 477 132 526 166
rect 560 132 576 166
rect 477 99 576 132
rect 612 166 944 183
rect 612 132 824 166
rect 858 132 944 166
rect 612 113 944 132
rect 119 73 441 79
rect 612 79 617 113
rect 651 79 689 113
rect 723 79 761 113
rect 795 79 833 113
rect 867 79 905 113
rect 939 79 944 113
rect 980 166 1030 221
rect 1014 132 1030 166
rect 980 99 1030 132
rect 612 73 944 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 140 701 174 735
rect 212 701 239 735
rect 239 701 246 735
rect 688 701 722 735
rect 760 701 794 735
rect 832 701 866 735
rect 904 701 938 735
rect 119 79 153 113
rect 191 79 225 113
rect 263 79 297 113
rect 335 79 369 113
rect 407 79 441 113
rect 617 79 651 113
rect 689 79 723 113
rect 761 79 795 113
rect 833 79 867 113
rect 905 79 939 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 735 1056 763
rect 0 701 140 735
rect 174 701 212 735
rect 246 701 688 735
rect 722 701 760 735
rect 794 701 832 735
rect 866 701 904 735
rect 938 701 1056 735
rect 0 689 1056 701
rect 0 113 1056 125
rect 0 79 119 113
rect 153 79 191 113
rect 225 79 263 113
rect 297 79 335 113
rect 369 79 407 113
rect 441 79 617 113
rect 651 79 689 113
rect 723 79 761 113
rect 795 79 833 113
rect 867 79 905 113
rect 939 79 1056 113
rect 0 51 1056 79
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2_1
flabel metal1 s 0 51 1056 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 1056 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 1056 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 1056 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 612 65 646 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1056 814
string GDS_END 249092
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 236720
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
