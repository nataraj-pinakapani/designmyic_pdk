magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< pwell >>
rect 10 66 1950 720
<< mvnmos >>
rect 228 92 328 694
rect 384 92 484 694
rect 540 92 640 694
rect 696 92 796 694
rect 852 92 952 694
rect 1008 92 1108 694
rect 1164 92 1264 694
rect 1320 92 1420 694
rect 1476 92 1576 694
rect 1632 92 1732 694
<< mvndiff >>
rect 172 682 228 694
rect 172 648 183 682
rect 217 648 228 682
rect 172 614 228 648
rect 172 580 183 614
rect 217 580 228 614
rect 172 546 228 580
rect 172 512 183 546
rect 217 512 228 546
rect 172 478 228 512
rect 172 444 183 478
rect 217 444 228 478
rect 172 410 228 444
rect 172 376 183 410
rect 217 376 228 410
rect 172 342 228 376
rect 172 308 183 342
rect 217 308 228 342
rect 172 274 228 308
rect 172 240 183 274
rect 217 240 228 274
rect 172 206 228 240
rect 172 172 183 206
rect 217 172 228 206
rect 172 138 228 172
rect 172 104 183 138
rect 217 104 228 138
rect 172 92 228 104
rect 328 682 384 694
rect 328 648 339 682
rect 373 648 384 682
rect 328 614 384 648
rect 328 580 339 614
rect 373 580 384 614
rect 328 546 384 580
rect 328 512 339 546
rect 373 512 384 546
rect 328 478 384 512
rect 328 444 339 478
rect 373 444 384 478
rect 328 410 384 444
rect 328 376 339 410
rect 373 376 384 410
rect 328 342 384 376
rect 328 308 339 342
rect 373 308 384 342
rect 328 274 384 308
rect 328 240 339 274
rect 373 240 384 274
rect 328 206 384 240
rect 328 172 339 206
rect 373 172 384 206
rect 328 138 384 172
rect 328 104 339 138
rect 373 104 384 138
rect 328 92 384 104
rect 484 682 540 694
rect 484 648 495 682
rect 529 648 540 682
rect 484 614 540 648
rect 484 580 495 614
rect 529 580 540 614
rect 484 546 540 580
rect 484 512 495 546
rect 529 512 540 546
rect 484 478 540 512
rect 484 444 495 478
rect 529 444 540 478
rect 484 410 540 444
rect 484 376 495 410
rect 529 376 540 410
rect 484 342 540 376
rect 484 308 495 342
rect 529 308 540 342
rect 484 274 540 308
rect 484 240 495 274
rect 529 240 540 274
rect 484 206 540 240
rect 484 172 495 206
rect 529 172 540 206
rect 484 138 540 172
rect 484 104 495 138
rect 529 104 540 138
rect 484 92 540 104
rect 640 682 696 694
rect 640 648 651 682
rect 685 648 696 682
rect 640 614 696 648
rect 640 580 651 614
rect 685 580 696 614
rect 640 546 696 580
rect 640 512 651 546
rect 685 512 696 546
rect 640 478 696 512
rect 640 444 651 478
rect 685 444 696 478
rect 640 410 696 444
rect 640 376 651 410
rect 685 376 696 410
rect 640 342 696 376
rect 640 308 651 342
rect 685 308 696 342
rect 640 274 696 308
rect 640 240 651 274
rect 685 240 696 274
rect 640 206 696 240
rect 640 172 651 206
rect 685 172 696 206
rect 640 138 696 172
rect 640 104 651 138
rect 685 104 696 138
rect 640 92 696 104
rect 796 682 852 694
rect 796 648 807 682
rect 841 648 852 682
rect 796 614 852 648
rect 796 580 807 614
rect 841 580 852 614
rect 796 546 852 580
rect 796 512 807 546
rect 841 512 852 546
rect 796 478 852 512
rect 796 444 807 478
rect 841 444 852 478
rect 796 410 852 444
rect 796 376 807 410
rect 841 376 852 410
rect 796 342 852 376
rect 796 308 807 342
rect 841 308 852 342
rect 796 274 852 308
rect 796 240 807 274
rect 841 240 852 274
rect 796 206 852 240
rect 796 172 807 206
rect 841 172 852 206
rect 796 138 852 172
rect 796 104 807 138
rect 841 104 852 138
rect 796 92 852 104
rect 952 682 1008 694
rect 952 648 963 682
rect 997 648 1008 682
rect 952 614 1008 648
rect 952 580 963 614
rect 997 580 1008 614
rect 952 546 1008 580
rect 952 512 963 546
rect 997 512 1008 546
rect 952 478 1008 512
rect 952 444 963 478
rect 997 444 1008 478
rect 952 410 1008 444
rect 952 376 963 410
rect 997 376 1008 410
rect 952 342 1008 376
rect 952 308 963 342
rect 997 308 1008 342
rect 952 274 1008 308
rect 952 240 963 274
rect 997 240 1008 274
rect 952 206 1008 240
rect 952 172 963 206
rect 997 172 1008 206
rect 952 138 1008 172
rect 952 104 963 138
rect 997 104 1008 138
rect 952 92 1008 104
rect 1108 682 1164 694
rect 1108 648 1119 682
rect 1153 648 1164 682
rect 1108 614 1164 648
rect 1108 580 1119 614
rect 1153 580 1164 614
rect 1108 546 1164 580
rect 1108 512 1119 546
rect 1153 512 1164 546
rect 1108 478 1164 512
rect 1108 444 1119 478
rect 1153 444 1164 478
rect 1108 410 1164 444
rect 1108 376 1119 410
rect 1153 376 1164 410
rect 1108 342 1164 376
rect 1108 308 1119 342
rect 1153 308 1164 342
rect 1108 274 1164 308
rect 1108 240 1119 274
rect 1153 240 1164 274
rect 1108 206 1164 240
rect 1108 172 1119 206
rect 1153 172 1164 206
rect 1108 138 1164 172
rect 1108 104 1119 138
rect 1153 104 1164 138
rect 1108 92 1164 104
rect 1264 682 1320 694
rect 1264 648 1275 682
rect 1309 648 1320 682
rect 1264 614 1320 648
rect 1264 580 1275 614
rect 1309 580 1320 614
rect 1264 546 1320 580
rect 1264 512 1275 546
rect 1309 512 1320 546
rect 1264 478 1320 512
rect 1264 444 1275 478
rect 1309 444 1320 478
rect 1264 410 1320 444
rect 1264 376 1275 410
rect 1309 376 1320 410
rect 1264 342 1320 376
rect 1264 308 1275 342
rect 1309 308 1320 342
rect 1264 274 1320 308
rect 1264 240 1275 274
rect 1309 240 1320 274
rect 1264 206 1320 240
rect 1264 172 1275 206
rect 1309 172 1320 206
rect 1264 138 1320 172
rect 1264 104 1275 138
rect 1309 104 1320 138
rect 1264 92 1320 104
rect 1420 682 1476 694
rect 1420 648 1431 682
rect 1465 648 1476 682
rect 1420 614 1476 648
rect 1420 580 1431 614
rect 1465 580 1476 614
rect 1420 546 1476 580
rect 1420 512 1431 546
rect 1465 512 1476 546
rect 1420 478 1476 512
rect 1420 444 1431 478
rect 1465 444 1476 478
rect 1420 410 1476 444
rect 1420 376 1431 410
rect 1465 376 1476 410
rect 1420 342 1476 376
rect 1420 308 1431 342
rect 1465 308 1476 342
rect 1420 274 1476 308
rect 1420 240 1431 274
rect 1465 240 1476 274
rect 1420 206 1476 240
rect 1420 172 1431 206
rect 1465 172 1476 206
rect 1420 138 1476 172
rect 1420 104 1431 138
rect 1465 104 1476 138
rect 1420 92 1476 104
rect 1576 682 1632 694
rect 1576 648 1587 682
rect 1621 648 1632 682
rect 1576 614 1632 648
rect 1576 580 1587 614
rect 1621 580 1632 614
rect 1576 546 1632 580
rect 1576 512 1587 546
rect 1621 512 1632 546
rect 1576 478 1632 512
rect 1576 444 1587 478
rect 1621 444 1632 478
rect 1576 410 1632 444
rect 1576 376 1587 410
rect 1621 376 1632 410
rect 1576 342 1632 376
rect 1576 308 1587 342
rect 1621 308 1632 342
rect 1576 274 1632 308
rect 1576 240 1587 274
rect 1621 240 1632 274
rect 1576 206 1632 240
rect 1576 172 1587 206
rect 1621 172 1632 206
rect 1576 138 1632 172
rect 1576 104 1587 138
rect 1621 104 1632 138
rect 1576 92 1632 104
rect 1732 682 1788 694
rect 1732 648 1743 682
rect 1777 648 1788 682
rect 1732 614 1788 648
rect 1732 580 1743 614
rect 1777 580 1788 614
rect 1732 546 1788 580
rect 1732 512 1743 546
rect 1777 512 1788 546
rect 1732 478 1788 512
rect 1732 444 1743 478
rect 1777 444 1788 478
rect 1732 410 1788 444
rect 1732 376 1743 410
rect 1777 376 1788 410
rect 1732 342 1788 376
rect 1732 308 1743 342
rect 1777 308 1788 342
rect 1732 274 1788 308
rect 1732 240 1743 274
rect 1777 240 1788 274
rect 1732 206 1788 240
rect 1732 172 1743 206
rect 1777 172 1788 206
rect 1732 138 1788 172
rect 1732 104 1743 138
rect 1777 104 1788 138
rect 1732 92 1788 104
<< mvndiffc >>
rect 183 648 217 682
rect 183 580 217 614
rect 183 512 217 546
rect 183 444 217 478
rect 183 376 217 410
rect 183 308 217 342
rect 183 240 217 274
rect 183 172 217 206
rect 183 104 217 138
rect 339 648 373 682
rect 339 580 373 614
rect 339 512 373 546
rect 339 444 373 478
rect 339 376 373 410
rect 339 308 373 342
rect 339 240 373 274
rect 339 172 373 206
rect 339 104 373 138
rect 495 648 529 682
rect 495 580 529 614
rect 495 512 529 546
rect 495 444 529 478
rect 495 376 529 410
rect 495 308 529 342
rect 495 240 529 274
rect 495 172 529 206
rect 495 104 529 138
rect 651 648 685 682
rect 651 580 685 614
rect 651 512 685 546
rect 651 444 685 478
rect 651 376 685 410
rect 651 308 685 342
rect 651 240 685 274
rect 651 172 685 206
rect 651 104 685 138
rect 807 648 841 682
rect 807 580 841 614
rect 807 512 841 546
rect 807 444 841 478
rect 807 376 841 410
rect 807 308 841 342
rect 807 240 841 274
rect 807 172 841 206
rect 807 104 841 138
rect 963 648 997 682
rect 963 580 997 614
rect 963 512 997 546
rect 963 444 997 478
rect 963 376 997 410
rect 963 308 997 342
rect 963 240 997 274
rect 963 172 997 206
rect 963 104 997 138
rect 1119 648 1153 682
rect 1119 580 1153 614
rect 1119 512 1153 546
rect 1119 444 1153 478
rect 1119 376 1153 410
rect 1119 308 1153 342
rect 1119 240 1153 274
rect 1119 172 1153 206
rect 1119 104 1153 138
rect 1275 648 1309 682
rect 1275 580 1309 614
rect 1275 512 1309 546
rect 1275 444 1309 478
rect 1275 376 1309 410
rect 1275 308 1309 342
rect 1275 240 1309 274
rect 1275 172 1309 206
rect 1275 104 1309 138
rect 1431 648 1465 682
rect 1431 580 1465 614
rect 1431 512 1465 546
rect 1431 444 1465 478
rect 1431 376 1465 410
rect 1431 308 1465 342
rect 1431 240 1465 274
rect 1431 172 1465 206
rect 1431 104 1465 138
rect 1587 648 1621 682
rect 1587 580 1621 614
rect 1587 512 1621 546
rect 1587 444 1621 478
rect 1587 376 1621 410
rect 1587 308 1621 342
rect 1587 240 1621 274
rect 1587 172 1621 206
rect 1587 104 1621 138
rect 1743 648 1777 682
rect 1743 580 1777 614
rect 1743 512 1777 546
rect 1743 444 1777 478
rect 1743 376 1777 410
rect 1743 308 1777 342
rect 1743 240 1777 274
rect 1743 172 1777 206
rect 1743 104 1777 138
<< mvpsubdiff >>
rect 36 648 94 694
rect 36 614 48 648
rect 82 614 94 648
rect 36 580 94 614
rect 36 546 48 580
rect 82 546 94 580
rect 36 512 94 546
rect 36 478 48 512
rect 82 478 94 512
rect 36 444 94 478
rect 36 410 48 444
rect 82 410 94 444
rect 36 376 94 410
rect 36 342 48 376
rect 82 342 94 376
rect 36 308 94 342
rect 36 274 48 308
rect 82 274 94 308
rect 36 240 94 274
rect 36 206 48 240
rect 82 206 94 240
rect 36 172 94 206
rect 36 138 48 172
rect 82 138 94 172
rect 36 92 94 138
rect 1866 648 1924 694
rect 1866 614 1878 648
rect 1912 614 1924 648
rect 1866 580 1924 614
rect 1866 546 1878 580
rect 1912 546 1924 580
rect 1866 512 1924 546
rect 1866 478 1878 512
rect 1912 478 1924 512
rect 1866 444 1924 478
rect 1866 410 1878 444
rect 1912 410 1924 444
rect 1866 376 1924 410
rect 1866 342 1878 376
rect 1912 342 1924 376
rect 1866 308 1924 342
rect 1866 274 1878 308
rect 1912 274 1924 308
rect 1866 240 1924 274
rect 1866 206 1878 240
rect 1912 206 1924 240
rect 1866 172 1924 206
rect 1866 138 1878 172
rect 1912 138 1924 172
rect 1866 92 1924 138
<< mvpsubdiffcont >>
rect 48 614 82 648
rect 48 546 82 580
rect 48 478 82 512
rect 48 410 82 444
rect 48 342 82 376
rect 48 274 82 308
rect 48 206 82 240
rect 48 138 82 172
rect 1878 614 1912 648
rect 1878 546 1912 580
rect 1878 478 1912 512
rect 1878 410 1912 444
rect 1878 342 1912 376
rect 1878 274 1912 308
rect 1878 206 1912 240
rect 1878 138 1912 172
<< poly >>
rect 199 766 1761 786
rect 199 732 215 766
rect 249 732 283 766
rect 317 732 351 766
rect 385 732 419 766
rect 453 732 487 766
rect 521 732 555 766
rect 589 732 623 766
rect 657 732 691 766
rect 725 732 759 766
rect 793 732 827 766
rect 861 732 895 766
rect 929 732 963 766
rect 997 732 1031 766
rect 1065 732 1099 766
rect 1133 732 1167 766
rect 1201 732 1235 766
rect 1269 732 1303 766
rect 1337 732 1371 766
rect 1405 732 1439 766
rect 1473 732 1507 766
rect 1541 732 1575 766
rect 1609 732 1643 766
rect 1677 732 1711 766
rect 1745 732 1761 766
rect 199 716 1761 732
rect 228 694 328 716
rect 384 694 484 716
rect 540 694 640 716
rect 696 694 796 716
rect 852 694 952 716
rect 1008 694 1108 716
rect 1164 694 1264 716
rect 1320 694 1420 716
rect 1476 694 1576 716
rect 1632 694 1732 716
rect 228 70 328 92
rect 384 70 484 92
rect 540 70 640 92
rect 696 70 796 92
rect 852 70 952 92
rect 1008 70 1108 92
rect 1164 70 1264 92
rect 1320 70 1420 92
rect 1476 70 1576 92
rect 1632 70 1732 92
rect 199 54 1761 70
rect 199 20 215 54
rect 249 20 283 54
rect 317 20 351 54
rect 385 20 419 54
rect 453 20 487 54
rect 521 20 555 54
rect 589 20 623 54
rect 657 20 691 54
rect 725 20 759 54
rect 793 20 827 54
rect 861 20 895 54
rect 929 20 963 54
rect 997 20 1031 54
rect 1065 20 1099 54
rect 1133 20 1167 54
rect 1201 20 1235 54
rect 1269 20 1303 54
rect 1337 20 1371 54
rect 1405 20 1439 54
rect 1473 20 1507 54
rect 1541 20 1575 54
rect 1609 20 1643 54
rect 1677 20 1711 54
rect 1745 20 1761 54
rect 199 0 1761 20
<< polycont >>
rect 215 732 249 766
rect 283 732 317 766
rect 351 732 385 766
rect 419 732 453 766
rect 487 732 521 766
rect 555 732 589 766
rect 623 732 657 766
rect 691 732 725 766
rect 759 732 793 766
rect 827 732 861 766
rect 895 732 929 766
rect 963 732 997 766
rect 1031 732 1065 766
rect 1099 732 1133 766
rect 1167 732 1201 766
rect 1235 732 1269 766
rect 1303 732 1337 766
rect 1371 732 1405 766
rect 1439 732 1473 766
rect 1507 732 1541 766
rect 1575 732 1609 766
rect 1643 732 1677 766
rect 1711 732 1745 766
rect 215 20 249 54
rect 283 20 317 54
rect 351 20 385 54
rect 419 20 453 54
rect 487 20 521 54
rect 555 20 589 54
rect 623 20 657 54
rect 691 20 725 54
rect 759 20 793 54
rect 827 20 861 54
rect 895 20 929 54
rect 963 20 997 54
rect 1031 20 1065 54
rect 1099 20 1133 54
rect 1167 20 1201 54
rect 1235 20 1269 54
rect 1303 20 1337 54
rect 1371 20 1405 54
rect 1439 20 1473 54
rect 1507 20 1541 54
rect 1575 20 1609 54
rect 1643 20 1677 54
rect 1711 20 1745 54
<< locali >>
rect 199 732 207 766
rect 249 732 279 766
rect 317 732 351 766
rect 385 732 419 766
rect 457 732 487 766
rect 529 732 555 766
rect 601 732 623 766
rect 673 732 691 766
rect 745 732 759 766
rect 817 732 827 766
rect 889 732 895 766
rect 961 732 963 766
rect 997 732 999 766
rect 1065 732 1071 766
rect 1133 732 1143 766
rect 1201 732 1215 766
rect 1269 732 1287 766
rect 1337 732 1359 766
rect 1405 732 1431 766
rect 1473 732 1503 766
rect 1541 732 1575 766
rect 1609 732 1643 766
rect 1681 732 1711 766
rect 1753 732 1761 766
rect 183 682 217 698
rect 48 662 82 664
rect 48 590 82 614
rect 48 518 82 546
rect 48 446 82 478
rect 48 376 82 410
rect 48 308 82 340
rect 48 240 82 268
rect 48 172 82 196
rect 48 122 82 124
rect 183 614 217 628
rect 183 546 217 556
rect 183 478 217 484
rect 183 410 217 412
rect 183 374 217 376
rect 183 302 217 308
rect 183 230 217 240
rect 183 158 217 172
rect 183 88 217 104
rect 339 682 373 698
rect 339 614 373 628
rect 339 546 373 556
rect 339 478 373 484
rect 339 410 373 412
rect 339 374 373 376
rect 339 302 373 308
rect 339 230 373 240
rect 339 158 373 172
rect 339 88 373 104
rect 495 682 529 698
rect 495 614 529 628
rect 495 546 529 556
rect 495 478 529 484
rect 495 410 529 412
rect 495 374 529 376
rect 495 302 529 308
rect 495 230 529 240
rect 495 158 529 172
rect 495 88 529 104
rect 651 682 685 698
rect 651 614 685 628
rect 651 546 685 556
rect 651 478 685 484
rect 651 410 685 412
rect 651 374 685 376
rect 651 302 685 308
rect 651 230 685 240
rect 651 158 685 172
rect 651 88 685 104
rect 807 682 841 698
rect 807 614 841 628
rect 807 546 841 556
rect 807 478 841 484
rect 807 410 841 412
rect 807 374 841 376
rect 807 302 841 308
rect 807 230 841 240
rect 807 158 841 172
rect 807 88 841 104
rect 963 682 997 698
rect 963 614 997 628
rect 963 546 997 556
rect 963 478 997 484
rect 963 410 997 412
rect 963 374 997 376
rect 963 302 997 308
rect 963 230 997 240
rect 963 158 997 172
rect 963 88 997 104
rect 1119 682 1153 698
rect 1119 614 1153 628
rect 1119 546 1153 556
rect 1119 478 1153 484
rect 1119 410 1153 412
rect 1119 374 1153 376
rect 1119 302 1153 308
rect 1119 230 1153 240
rect 1119 158 1153 172
rect 1119 88 1153 104
rect 1275 682 1309 698
rect 1275 614 1309 628
rect 1275 546 1309 556
rect 1275 478 1309 484
rect 1275 410 1309 412
rect 1275 374 1309 376
rect 1275 302 1309 308
rect 1275 230 1309 240
rect 1275 158 1309 172
rect 1275 88 1309 104
rect 1431 682 1465 698
rect 1431 614 1465 628
rect 1431 546 1465 556
rect 1431 478 1465 484
rect 1431 410 1465 412
rect 1431 374 1465 376
rect 1431 302 1465 308
rect 1431 230 1465 240
rect 1431 158 1465 172
rect 1431 88 1465 104
rect 1587 682 1621 698
rect 1587 614 1621 628
rect 1587 546 1621 556
rect 1587 478 1621 484
rect 1587 410 1621 412
rect 1587 374 1621 376
rect 1587 302 1621 308
rect 1587 230 1621 240
rect 1587 158 1621 172
rect 1587 88 1621 104
rect 1743 682 1777 698
rect 1743 614 1777 628
rect 1743 546 1777 556
rect 1743 478 1777 484
rect 1743 410 1777 412
rect 1743 374 1777 376
rect 1743 302 1777 308
rect 1743 230 1777 240
rect 1743 158 1777 172
rect 1878 662 1912 664
rect 1878 590 1912 614
rect 1878 518 1912 546
rect 1878 446 1912 478
rect 1878 376 1912 410
rect 1878 308 1912 340
rect 1878 240 1912 268
rect 1878 172 1912 196
rect 1878 122 1912 124
rect 1743 88 1777 104
rect 199 20 207 54
rect 249 20 279 54
rect 317 20 351 54
rect 385 20 419 54
rect 457 20 487 54
rect 529 20 555 54
rect 601 20 623 54
rect 673 20 691 54
rect 745 20 759 54
rect 817 20 827 54
rect 889 20 895 54
rect 961 20 963 54
rect 997 20 999 54
rect 1065 20 1071 54
rect 1133 20 1143 54
rect 1201 20 1215 54
rect 1269 20 1287 54
rect 1337 20 1359 54
rect 1405 20 1431 54
rect 1473 20 1503 54
rect 1541 20 1575 54
rect 1609 20 1643 54
rect 1681 20 1711 54
rect 1753 20 1761 54
<< viali >>
rect 207 732 215 766
rect 215 732 241 766
rect 279 732 283 766
rect 283 732 313 766
rect 351 732 385 766
rect 423 732 453 766
rect 453 732 457 766
rect 495 732 521 766
rect 521 732 529 766
rect 567 732 589 766
rect 589 732 601 766
rect 639 732 657 766
rect 657 732 673 766
rect 711 732 725 766
rect 725 732 745 766
rect 783 732 793 766
rect 793 732 817 766
rect 855 732 861 766
rect 861 732 889 766
rect 927 732 929 766
rect 929 732 961 766
rect 999 732 1031 766
rect 1031 732 1033 766
rect 1071 732 1099 766
rect 1099 732 1105 766
rect 1143 732 1167 766
rect 1167 732 1177 766
rect 1215 732 1235 766
rect 1235 732 1249 766
rect 1287 732 1303 766
rect 1303 732 1321 766
rect 1359 732 1371 766
rect 1371 732 1393 766
rect 1431 732 1439 766
rect 1439 732 1465 766
rect 1503 732 1507 766
rect 1507 732 1537 766
rect 1575 732 1609 766
rect 1647 732 1677 766
rect 1677 732 1681 766
rect 1719 732 1745 766
rect 1745 732 1753 766
rect 48 648 82 662
rect 48 628 82 648
rect 48 580 82 590
rect 48 556 82 580
rect 48 512 82 518
rect 48 484 82 512
rect 48 444 82 446
rect 48 412 82 444
rect 48 342 82 374
rect 48 340 82 342
rect 48 274 82 302
rect 48 268 82 274
rect 48 206 82 230
rect 48 196 82 206
rect 48 138 82 158
rect 48 124 82 138
rect 183 648 217 662
rect 183 628 217 648
rect 183 580 217 590
rect 183 556 217 580
rect 183 512 217 518
rect 183 484 217 512
rect 183 444 217 446
rect 183 412 217 444
rect 183 342 217 374
rect 183 340 217 342
rect 183 274 217 302
rect 183 268 217 274
rect 183 206 217 230
rect 183 196 217 206
rect 183 138 217 158
rect 183 124 217 138
rect 339 648 373 662
rect 339 628 373 648
rect 339 580 373 590
rect 339 556 373 580
rect 339 512 373 518
rect 339 484 373 512
rect 339 444 373 446
rect 339 412 373 444
rect 339 342 373 374
rect 339 340 373 342
rect 339 274 373 302
rect 339 268 373 274
rect 339 206 373 230
rect 339 196 373 206
rect 339 138 373 158
rect 339 124 373 138
rect 495 648 529 662
rect 495 628 529 648
rect 495 580 529 590
rect 495 556 529 580
rect 495 512 529 518
rect 495 484 529 512
rect 495 444 529 446
rect 495 412 529 444
rect 495 342 529 374
rect 495 340 529 342
rect 495 274 529 302
rect 495 268 529 274
rect 495 206 529 230
rect 495 196 529 206
rect 495 138 529 158
rect 495 124 529 138
rect 651 648 685 662
rect 651 628 685 648
rect 651 580 685 590
rect 651 556 685 580
rect 651 512 685 518
rect 651 484 685 512
rect 651 444 685 446
rect 651 412 685 444
rect 651 342 685 374
rect 651 340 685 342
rect 651 274 685 302
rect 651 268 685 274
rect 651 206 685 230
rect 651 196 685 206
rect 651 138 685 158
rect 651 124 685 138
rect 807 648 841 662
rect 807 628 841 648
rect 807 580 841 590
rect 807 556 841 580
rect 807 512 841 518
rect 807 484 841 512
rect 807 444 841 446
rect 807 412 841 444
rect 807 342 841 374
rect 807 340 841 342
rect 807 274 841 302
rect 807 268 841 274
rect 807 206 841 230
rect 807 196 841 206
rect 807 138 841 158
rect 807 124 841 138
rect 963 648 997 662
rect 963 628 997 648
rect 963 580 997 590
rect 963 556 997 580
rect 963 512 997 518
rect 963 484 997 512
rect 963 444 997 446
rect 963 412 997 444
rect 963 342 997 374
rect 963 340 997 342
rect 963 274 997 302
rect 963 268 997 274
rect 963 206 997 230
rect 963 196 997 206
rect 963 138 997 158
rect 963 124 997 138
rect 1119 648 1153 662
rect 1119 628 1153 648
rect 1119 580 1153 590
rect 1119 556 1153 580
rect 1119 512 1153 518
rect 1119 484 1153 512
rect 1119 444 1153 446
rect 1119 412 1153 444
rect 1119 342 1153 374
rect 1119 340 1153 342
rect 1119 274 1153 302
rect 1119 268 1153 274
rect 1119 206 1153 230
rect 1119 196 1153 206
rect 1119 138 1153 158
rect 1119 124 1153 138
rect 1275 648 1309 662
rect 1275 628 1309 648
rect 1275 580 1309 590
rect 1275 556 1309 580
rect 1275 512 1309 518
rect 1275 484 1309 512
rect 1275 444 1309 446
rect 1275 412 1309 444
rect 1275 342 1309 374
rect 1275 340 1309 342
rect 1275 274 1309 302
rect 1275 268 1309 274
rect 1275 206 1309 230
rect 1275 196 1309 206
rect 1275 138 1309 158
rect 1275 124 1309 138
rect 1431 648 1465 662
rect 1431 628 1465 648
rect 1431 580 1465 590
rect 1431 556 1465 580
rect 1431 512 1465 518
rect 1431 484 1465 512
rect 1431 444 1465 446
rect 1431 412 1465 444
rect 1431 342 1465 374
rect 1431 340 1465 342
rect 1431 274 1465 302
rect 1431 268 1465 274
rect 1431 206 1465 230
rect 1431 196 1465 206
rect 1431 138 1465 158
rect 1431 124 1465 138
rect 1587 648 1621 662
rect 1587 628 1621 648
rect 1587 580 1621 590
rect 1587 556 1621 580
rect 1587 512 1621 518
rect 1587 484 1621 512
rect 1587 444 1621 446
rect 1587 412 1621 444
rect 1587 342 1621 374
rect 1587 340 1621 342
rect 1587 274 1621 302
rect 1587 268 1621 274
rect 1587 206 1621 230
rect 1587 196 1621 206
rect 1587 138 1621 158
rect 1587 124 1621 138
rect 1743 648 1777 662
rect 1743 628 1777 648
rect 1743 580 1777 590
rect 1743 556 1777 580
rect 1743 512 1777 518
rect 1743 484 1777 512
rect 1743 444 1777 446
rect 1743 412 1777 444
rect 1743 342 1777 374
rect 1743 340 1777 342
rect 1743 274 1777 302
rect 1743 268 1777 274
rect 1743 206 1777 230
rect 1743 196 1777 206
rect 1743 138 1777 158
rect 1743 124 1777 138
rect 1878 648 1912 662
rect 1878 628 1912 648
rect 1878 580 1912 590
rect 1878 556 1912 580
rect 1878 512 1912 518
rect 1878 484 1912 512
rect 1878 444 1912 446
rect 1878 412 1912 444
rect 1878 342 1912 374
rect 1878 340 1912 342
rect 1878 274 1912 302
rect 1878 268 1912 274
rect 1878 206 1912 230
rect 1878 196 1912 206
rect 1878 138 1912 158
rect 1878 124 1912 138
rect 207 20 215 54
rect 215 20 241 54
rect 279 20 283 54
rect 283 20 313 54
rect 351 20 385 54
rect 423 20 453 54
rect 453 20 457 54
rect 495 20 521 54
rect 521 20 529 54
rect 567 20 589 54
rect 589 20 601 54
rect 639 20 657 54
rect 657 20 673 54
rect 711 20 725 54
rect 725 20 745 54
rect 783 20 793 54
rect 793 20 817 54
rect 855 20 861 54
rect 861 20 889 54
rect 927 20 929 54
rect 929 20 961 54
rect 999 20 1031 54
rect 1031 20 1033 54
rect 1071 20 1099 54
rect 1099 20 1105 54
rect 1143 20 1167 54
rect 1167 20 1177 54
rect 1215 20 1235 54
rect 1235 20 1249 54
rect 1287 20 1303 54
rect 1303 20 1321 54
rect 1359 20 1371 54
rect 1371 20 1393 54
rect 1431 20 1439 54
rect 1439 20 1465 54
rect 1503 20 1507 54
rect 1507 20 1537 54
rect 1575 20 1609 54
rect 1647 20 1677 54
rect 1677 20 1681 54
rect 1719 20 1745 54
rect 1745 20 1753 54
<< metal1 >>
rect 195 766 1765 786
rect 195 732 207 766
rect 241 732 279 766
rect 313 732 351 766
rect 385 732 423 766
rect 457 732 495 766
rect 529 732 567 766
rect 601 732 639 766
rect 673 732 711 766
rect 745 732 783 766
rect 817 732 855 766
rect 889 732 927 766
rect 961 732 999 766
rect 1033 732 1071 766
rect 1105 732 1143 766
rect 1177 732 1215 766
rect 1249 732 1287 766
rect 1321 732 1359 766
rect 1393 732 1431 766
rect 1465 732 1503 766
rect 1537 732 1575 766
rect 1609 732 1647 766
rect 1681 732 1719 766
rect 1753 732 1765 766
rect 195 720 1765 732
rect 36 662 94 674
rect 36 628 48 662
rect 82 628 94 662
rect 36 590 94 628
rect 36 556 48 590
rect 82 556 94 590
rect 36 518 94 556
rect 36 484 48 518
rect 82 484 94 518
rect 36 446 94 484
rect 36 412 48 446
rect 82 412 94 446
rect 36 374 94 412
rect 36 340 48 374
rect 82 340 94 374
rect 36 302 94 340
rect 36 268 48 302
rect 82 268 94 302
rect 36 230 94 268
rect 36 196 48 230
rect 82 196 94 230
rect 36 158 94 196
rect 36 124 48 158
rect 82 124 94 158
rect 36 112 94 124
rect 174 662 226 674
rect 174 628 183 662
rect 217 628 226 662
rect 174 590 226 628
rect 174 556 183 590
rect 217 556 226 590
rect 174 518 226 556
rect 174 484 183 518
rect 217 484 226 518
rect 174 446 226 484
rect 174 412 183 446
rect 217 412 226 446
rect 174 374 226 412
rect 174 362 183 374
rect 217 362 226 374
rect 174 302 226 310
rect 174 298 183 302
rect 217 298 226 302
rect 174 234 226 246
rect 174 170 226 182
rect 174 112 226 118
rect 330 668 382 674
rect 330 604 382 616
rect 330 540 382 552
rect 330 484 339 488
rect 373 484 382 488
rect 330 476 382 484
rect 330 412 339 424
rect 373 412 382 424
rect 330 374 382 412
rect 330 340 339 374
rect 373 340 382 374
rect 330 302 382 340
rect 330 268 339 302
rect 373 268 382 302
rect 330 230 382 268
rect 330 196 339 230
rect 373 196 382 230
rect 330 158 382 196
rect 330 124 339 158
rect 373 124 382 158
rect 330 112 382 124
rect 486 662 538 674
rect 486 628 495 662
rect 529 628 538 662
rect 486 590 538 628
rect 486 556 495 590
rect 529 556 538 590
rect 486 518 538 556
rect 486 484 495 518
rect 529 484 538 518
rect 486 446 538 484
rect 486 412 495 446
rect 529 412 538 446
rect 486 374 538 412
rect 486 362 495 374
rect 529 362 538 374
rect 486 302 538 310
rect 486 298 495 302
rect 529 298 538 302
rect 486 234 538 246
rect 486 170 538 182
rect 486 112 538 118
rect 642 668 694 674
rect 642 604 694 616
rect 642 540 694 552
rect 642 484 651 488
rect 685 484 694 488
rect 642 476 694 484
rect 642 412 651 424
rect 685 412 694 424
rect 642 374 694 412
rect 642 340 651 374
rect 685 340 694 374
rect 642 302 694 340
rect 642 268 651 302
rect 685 268 694 302
rect 642 230 694 268
rect 642 196 651 230
rect 685 196 694 230
rect 642 158 694 196
rect 642 124 651 158
rect 685 124 694 158
rect 642 112 694 124
rect 798 662 850 674
rect 798 628 807 662
rect 841 628 850 662
rect 798 590 850 628
rect 798 556 807 590
rect 841 556 850 590
rect 798 518 850 556
rect 798 484 807 518
rect 841 484 850 518
rect 798 446 850 484
rect 798 412 807 446
rect 841 412 850 446
rect 798 374 850 412
rect 798 362 807 374
rect 841 362 850 374
rect 798 302 850 310
rect 798 298 807 302
rect 841 298 850 302
rect 798 234 850 246
rect 798 170 850 182
rect 798 112 850 118
rect 954 668 1006 674
rect 954 604 1006 616
rect 954 540 1006 552
rect 954 484 963 488
rect 997 484 1006 488
rect 954 476 1006 484
rect 954 412 963 424
rect 997 412 1006 424
rect 954 374 1006 412
rect 954 340 963 374
rect 997 340 1006 374
rect 954 302 1006 340
rect 954 268 963 302
rect 997 268 1006 302
rect 954 230 1006 268
rect 954 196 963 230
rect 997 196 1006 230
rect 954 158 1006 196
rect 954 124 963 158
rect 997 124 1006 158
rect 954 112 1006 124
rect 1110 662 1162 674
rect 1110 628 1119 662
rect 1153 628 1162 662
rect 1110 590 1162 628
rect 1110 556 1119 590
rect 1153 556 1162 590
rect 1110 518 1162 556
rect 1110 484 1119 518
rect 1153 484 1162 518
rect 1110 446 1162 484
rect 1110 412 1119 446
rect 1153 412 1162 446
rect 1110 374 1162 412
rect 1110 362 1119 374
rect 1153 362 1162 374
rect 1110 302 1162 310
rect 1110 298 1119 302
rect 1153 298 1162 302
rect 1110 234 1162 246
rect 1110 170 1162 182
rect 1110 112 1162 118
rect 1266 668 1318 674
rect 1266 604 1318 616
rect 1266 540 1318 552
rect 1266 484 1275 488
rect 1309 484 1318 488
rect 1266 476 1318 484
rect 1266 412 1275 424
rect 1309 412 1318 424
rect 1266 374 1318 412
rect 1266 340 1275 374
rect 1309 340 1318 374
rect 1266 302 1318 340
rect 1266 268 1275 302
rect 1309 268 1318 302
rect 1266 230 1318 268
rect 1266 196 1275 230
rect 1309 196 1318 230
rect 1266 158 1318 196
rect 1266 124 1275 158
rect 1309 124 1318 158
rect 1266 112 1318 124
rect 1422 662 1474 674
rect 1422 628 1431 662
rect 1465 628 1474 662
rect 1422 590 1474 628
rect 1422 556 1431 590
rect 1465 556 1474 590
rect 1422 518 1474 556
rect 1422 484 1431 518
rect 1465 484 1474 518
rect 1422 446 1474 484
rect 1422 412 1431 446
rect 1465 412 1474 446
rect 1422 374 1474 412
rect 1422 362 1431 374
rect 1465 362 1474 374
rect 1422 302 1474 310
rect 1422 298 1431 302
rect 1465 298 1474 302
rect 1422 234 1474 246
rect 1422 170 1474 182
rect 1422 112 1474 118
rect 1578 668 1630 674
rect 1578 604 1630 616
rect 1578 540 1630 552
rect 1578 484 1587 488
rect 1621 484 1630 488
rect 1578 476 1630 484
rect 1578 412 1587 424
rect 1621 412 1630 424
rect 1578 374 1630 412
rect 1578 340 1587 374
rect 1621 340 1630 374
rect 1578 302 1630 340
rect 1578 268 1587 302
rect 1621 268 1630 302
rect 1578 230 1630 268
rect 1578 196 1587 230
rect 1621 196 1630 230
rect 1578 158 1630 196
rect 1578 124 1587 158
rect 1621 124 1630 158
rect 1578 112 1630 124
rect 1734 662 1786 674
rect 1734 628 1743 662
rect 1777 628 1786 662
rect 1734 590 1786 628
rect 1734 556 1743 590
rect 1777 556 1786 590
rect 1734 518 1786 556
rect 1734 484 1743 518
rect 1777 484 1786 518
rect 1734 446 1786 484
rect 1734 412 1743 446
rect 1777 412 1786 446
rect 1734 374 1786 412
rect 1734 362 1743 374
rect 1777 362 1786 374
rect 1734 302 1786 310
rect 1734 298 1743 302
rect 1777 298 1786 302
rect 1734 234 1786 246
rect 1734 170 1786 182
rect 1734 112 1786 118
rect 1866 662 1924 674
rect 1866 628 1878 662
rect 1912 628 1924 662
rect 1866 590 1924 628
rect 1866 556 1878 590
rect 1912 556 1924 590
rect 1866 518 1924 556
rect 1866 484 1878 518
rect 1912 484 1924 518
rect 1866 446 1924 484
rect 1866 412 1878 446
rect 1912 412 1924 446
rect 1866 374 1924 412
rect 1866 340 1878 374
rect 1912 340 1924 374
rect 1866 302 1924 340
rect 1866 268 1878 302
rect 1912 268 1924 302
rect 1866 230 1924 268
rect 1866 196 1878 230
rect 1912 196 1924 230
rect 1866 158 1924 196
rect 1866 124 1878 158
rect 1912 124 1924 158
rect 1866 112 1924 124
rect 195 54 1765 66
rect 195 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1765 54
rect 195 0 1765 20
<< via1 >>
rect 174 340 183 362
rect 183 340 217 362
rect 217 340 226 362
rect 174 310 226 340
rect 174 268 183 298
rect 183 268 217 298
rect 217 268 226 298
rect 174 246 226 268
rect 174 230 226 234
rect 174 196 183 230
rect 183 196 217 230
rect 217 196 226 230
rect 174 182 226 196
rect 174 158 226 170
rect 174 124 183 158
rect 183 124 217 158
rect 217 124 226 158
rect 174 118 226 124
rect 330 662 382 668
rect 330 628 339 662
rect 339 628 373 662
rect 373 628 382 662
rect 330 616 382 628
rect 330 590 382 604
rect 330 556 339 590
rect 339 556 373 590
rect 373 556 382 590
rect 330 552 382 556
rect 330 518 382 540
rect 330 488 339 518
rect 339 488 373 518
rect 373 488 382 518
rect 330 446 382 476
rect 330 424 339 446
rect 339 424 373 446
rect 373 424 382 446
rect 486 340 495 362
rect 495 340 529 362
rect 529 340 538 362
rect 486 310 538 340
rect 486 268 495 298
rect 495 268 529 298
rect 529 268 538 298
rect 486 246 538 268
rect 486 230 538 234
rect 486 196 495 230
rect 495 196 529 230
rect 529 196 538 230
rect 486 182 538 196
rect 486 158 538 170
rect 486 124 495 158
rect 495 124 529 158
rect 529 124 538 158
rect 486 118 538 124
rect 642 662 694 668
rect 642 628 651 662
rect 651 628 685 662
rect 685 628 694 662
rect 642 616 694 628
rect 642 590 694 604
rect 642 556 651 590
rect 651 556 685 590
rect 685 556 694 590
rect 642 552 694 556
rect 642 518 694 540
rect 642 488 651 518
rect 651 488 685 518
rect 685 488 694 518
rect 642 446 694 476
rect 642 424 651 446
rect 651 424 685 446
rect 685 424 694 446
rect 798 340 807 362
rect 807 340 841 362
rect 841 340 850 362
rect 798 310 850 340
rect 798 268 807 298
rect 807 268 841 298
rect 841 268 850 298
rect 798 246 850 268
rect 798 230 850 234
rect 798 196 807 230
rect 807 196 841 230
rect 841 196 850 230
rect 798 182 850 196
rect 798 158 850 170
rect 798 124 807 158
rect 807 124 841 158
rect 841 124 850 158
rect 798 118 850 124
rect 954 662 1006 668
rect 954 628 963 662
rect 963 628 997 662
rect 997 628 1006 662
rect 954 616 1006 628
rect 954 590 1006 604
rect 954 556 963 590
rect 963 556 997 590
rect 997 556 1006 590
rect 954 552 1006 556
rect 954 518 1006 540
rect 954 488 963 518
rect 963 488 997 518
rect 997 488 1006 518
rect 954 446 1006 476
rect 954 424 963 446
rect 963 424 997 446
rect 997 424 1006 446
rect 1110 340 1119 362
rect 1119 340 1153 362
rect 1153 340 1162 362
rect 1110 310 1162 340
rect 1110 268 1119 298
rect 1119 268 1153 298
rect 1153 268 1162 298
rect 1110 246 1162 268
rect 1110 230 1162 234
rect 1110 196 1119 230
rect 1119 196 1153 230
rect 1153 196 1162 230
rect 1110 182 1162 196
rect 1110 158 1162 170
rect 1110 124 1119 158
rect 1119 124 1153 158
rect 1153 124 1162 158
rect 1110 118 1162 124
rect 1266 662 1318 668
rect 1266 628 1275 662
rect 1275 628 1309 662
rect 1309 628 1318 662
rect 1266 616 1318 628
rect 1266 590 1318 604
rect 1266 556 1275 590
rect 1275 556 1309 590
rect 1309 556 1318 590
rect 1266 552 1318 556
rect 1266 518 1318 540
rect 1266 488 1275 518
rect 1275 488 1309 518
rect 1309 488 1318 518
rect 1266 446 1318 476
rect 1266 424 1275 446
rect 1275 424 1309 446
rect 1309 424 1318 446
rect 1422 340 1431 362
rect 1431 340 1465 362
rect 1465 340 1474 362
rect 1422 310 1474 340
rect 1422 268 1431 298
rect 1431 268 1465 298
rect 1465 268 1474 298
rect 1422 246 1474 268
rect 1422 230 1474 234
rect 1422 196 1431 230
rect 1431 196 1465 230
rect 1465 196 1474 230
rect 1422 182 1474 196
rect 1422 158 1474 170
rect 1422 124 1431 158
rect 1431 124 1465 158
rect 1465 124 1474 158
rect 1422 118 1474 124
rect 1578 662 1630 668
rect 1578 628 1587 662
rect 1587 628 1621 662
rect 1621 628 1630 662
rect 1578 616 1630 628
rect 1578 590 1630 604
rect 1578 556 1587 590
rect 1587 556 1621 590
rect 1621 556 1630 590
rect 1578 552 1630 556
rect 1578 518 1630 540
rect 1578 488 1587 518
rect 1587 488 1621 518
rect 1621 488 1630 518
rect 1578 446 1630 476
rect 1578 424 1587 446
rect 1587 424 1621 446
rect 1621 424 1630 446
rect 1734 340 1743 362
rect 1743 340 1777 362
rect 1777 340 1786 362
rect 1734 310 1786 340
rect 1734 268 1743 298
rect 1743 268 1777 298
rect 1777 268 1786 298
rect 1734 246 1786 268
rect 1734 230 1786 234
rect 1734 196 1743 230
rect 1743 196 1777 230
rect 1777 196 1786 230
rect 1734 182 1786 196
rect 1734 158 1786 170
rect 1734 124 1743 158
rect 1743 124 1777 158
rect 1777 124 1786 158
rect 1734 118 1786 124
<< metal2 >>
rect 10 668 1950 674
rect 10 616 330 668
rect 382 616 642 668
rect 694 616 954 668
rect 1006 616 1266 668
rect 1318 616 1578 668
rect 1630 616 1950 668
rect 10 604 1950 616
rect 10 552 330 604
rect 382 552 642 604
rect 694 552 954 604
rect 1006 552 1266 604
rect 1318 552 1578 604
rect 1630 552 1950 604
rect 10 540 1950 552
rect 10 488 330 540
rect 382 488 642 540
rect 694 488 954 540
rect 1006 488 1266 540
rect 1318 488 1578 540
rect 1630 488 1950 540
rect 10 476 1950 488
rect 10 424 330 476
rect 382 424 642 476
rect 694 424 954 476
rect 1006 424 1266 476
rect 1318 424 1578 476
rect 1630 424 1950 476
rect 10 418 1950 424
rect 10 362 1950 368
rect 10 310 174 362
rect 226 310 486 362
rect 538 310 798 362
rect 850 310 1110 362
rect 1162 310 1422 362
rect 1474 310 1734 362
rect 1786 310 1950 362
rect 10 298 1950 310
rect 10 246 174 298
rect 226 246 486 298
rect 538 246 798 298
rect 850 246 1110 298
rect 1162 246 1422 298
rect 1474 246 1734 298
rect 1786 246 1950 298
rect 10 234 1950 246
rect 10 182 174 234
rect 226 182 486 234
rect 538 182 798 234
rect 850 182 1110 234
rect 1162 182 1422 234
rect 1474 182 1734 234
rect 1786 182 1950 234
rect 10 170 1950 182
rect 10 118 174 170
rect 226 118 486 170
rect 538 118 798 170
rect 850 118 1110 170
rect 1162 118 1422 170
rect 1474 118 1734 170
rect 1786 118 1950 170
rect 10 112 1950 118
<< labels >>
flabel comment s 356 393 356 393 0 FreeSans 300 0 0 0 D
flabel comment s 356 393 356 393 0 FreeSans 300 0 0 0 S
flabel comment s 200 393 200 393 0 FreeSans 300 0 0 0 S
flabel comment s 200 393 200 393 0 FreeSans 300 0 0 0 S
flabel comment s 668 393 668 393 0 FreeSans 300 0 0 0 D
flabel comment s 512 393 512 393 0 FreeSans 300 0 0 0 S
flabel comment s 668 393 668 393 0 FreeSans 300 0 0 0 S
flabel comment s 512 393 512 393 0 FreeSans 300 0 0 0 S
flabel comment s 1136 393 1136 393 0 FreeSans 300 0 0 0 D
flabel comment s 980 393 980 393 0 FreeSans 300 0 0 0 S
flabel comment s 824 393 824 393 0 FreeSans 300 0 0 0 D
flabel comment s 1136 393 1136 393 0 FreeSans 300 0 0 0 S
flabel comment s 980 393 980 393 0 FreeSans 300 0 0 0 S
flabel comment s 824 393 824 393 0 FreeSans 300 0 0 0 S
flabel comment s 1292 393 1292 393 0 FreeSans 300 0 0 0 S
flabel comment s 1448 393 1448 393 0 FreeSans 300 0 0 0 S
flabel comment s 1604 393 1604 393 0 FreeSans 300 0 0 0 S
flabel comment s 1292 393 1292 393 0 FreeSans 300 0 0 0 D
flabel comment s 1448 393 1448 393 0 FreeSans 300 0 0 0 S
flabel comment s 1604 393 1604 393 0 FreeSans 300 0 0 0 D
flabel comment s 1760 393 1760 393 0 FreeSans 300 0 0 0 S
flabel metal2 s 31 219 142 267 0 FreeSans 200 0 0 0 SOURCE
port 1 nsew
flabel metal2 s 28 514 125 567 0 FreeSans 200 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 1884 318 1914 468 0 FreeSans 200 90 0 0 SUBSTRATE
port 3 nsew
flabel metal1 s 927 734 1049 767 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 929 14 1026 49 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 56 326 82 455 0 FreeSans 200 90 0 0 SUBSTRATE
port 3 nsew
<< properties >>
string GDS_END 4379702
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_pr/sky130_fd_pr.gds
string GDS_START 4348248
<< end >>
