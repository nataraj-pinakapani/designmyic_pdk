magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 21 799 731 1967
<< pwell >>
rect 81 76 535 728
<< mvnmos >>
rect 160 102 280 702
rect 336 102 456 702
<< mvpmos >>
rect 140 865 260 1865
rect 316 865 436 1865
rect 492 865 612 1865
<< mvndiff >>
rect 107 624 160 702
rect 107 590 115 624
rect 149 590 160 624
rect 107 556 160 590
rect 107 522 115 556
rect 149 522 160 556
rect 107 488 160 522
rect 107 454 115 488
rect 149 454 160 488
rect 107 420 160 454
rect 107 386 115 420
rect 149 386 160 420
rect 107 352 160 386
rect 107 318 115 352
rect 149 318 160 352
rect 107 284 160 318
rect 107 250 115 284
rect 149 250 160 284
rect 107 216 160 250
rect 107 182 115 216
rect 149 182 160 216
rect 107 148 160 182
rect 107 114 115 148
rect 149 114 160 148
rect 107 102 160 114
rect 280 624 336 702
rect 280 590 291 624
rect 325 590 336 624
rect 280 556 336 590
rect 280 522 291 556
rect 325 522 336 556
rect 280 488 336 522
rect 280 454 291 488
rect 325 454 336 488
rect 280 420 336 454
rect 280 386 291 420
rect 325 386 336 420
rect 280 352 336 386
rect 280 318 291 352
rect 325 318 336 352
rect 280 284 336 318
rect 280 250 291 284
rect 325 250 336 284
rect 280 216 336 250
rect 280 182 291 216
rect 325 182 336 216
rect 280 148 336 182
rect 280 114 291 148
rect 325 114 336 148
rect 280 102 336 114
rect 456 624 509 702
rect 456 590 467 624
rect 501 590 509 624
rect 456 556 509 590
rect 456 522 467 556
rect 501 522 509 556
rect 456 488 509 522
rect 456 454 467 488
rect 501 454 509 488
rect 456 420 509 454
rect 456 386 467 420
rect 501 386 509 420
rect 456 352 509 386
rect 456 318 467 352
rect 501 318 509 352
rect 456 284 509 318
rect 456 250 467 284
rect 501 250 509 284
rect 456 216 509 250
rect 456 182 467 216
rect 501 182 509 216
rect 456 148 509 182
rect 456 114 467 148
rect 501 114 509 148
rect 456 102 509 114
<< mvpdiff >>
rect 87 1853 140 1865
rect 87 1819 95 1853
rect 129 1819 140 1853
rect 87 1785 140 1819
rect 87 1751 95 1785
rect 129 1751 140 1785
rect 87 1717 140 1751
rect 87 1683 95 1717
rect 129 1683 140 1717
rect 87 1649 140 1683
rect 87 1615 95 1649
rect 129 1615 140 1649
rect 87 1581 140 1615
rect 87 1547 95 1581
rect 129 1547 140 1581
rect 87 1513 140 1547
rect 87 1479 95 1513
rect 129 1479 140 1513
rect 87 1445 140 1479
rect 87 1411 95 1445
rect 129 1411 140 1445
rect 87 1377 140 1411
rect 87 1343 95 1377
rect 129 1343 140 1377
rect 87 1309 140 1343
rect 87 1275 95 1309
rect 129 1275 140 1309
rect 87 1241 140 1275
rect 87 1207 95 1241
rect 129 1207 140 1241
rect 87 1173 140 1207
rect 87 1139 95 1173
rect 129 1139 140 1173
rect 87 1105 140 1139
rect 87 1071 95 1105
rect 129 1071 140 1105
rect 87 1037 140 1071
rect 87 1003 95 1037
rect 129 1003 140 1037
rect 87 969 140 1003
rect 87 935 95 969
rect 129 935 140 969
rect 87 865 140 935
rect 260 1853 316 1865
rect 260 1819 271 1853
rect 305 1819 316 1853
rect 260 1785 316 1819
rect 260 1751 271 1785
rect 305 1751 316 1785
rect 260 1717 316 1751
rect 260 1683 271 1717
rect 305 1683 316 1717
rect 260 1649 316 1683
rect 260 1615 271 1649
rect 305 1615 316 1649
rect 260 1581 316 1615
rect 260 1547 271 1581
rect 305 1547 316 1581
rect 260 1513 316 1547
rect 260 1479 271 1513
rect 305 1479 316 1513
rect 260 1445 316 1479
rect 260 1411 271 1445
rect 305 1411 316 1445
rect 260 1377 316 1411
rect 260 1343 271 1377
rect 305 1343 316 1377
rect 260 1309 316 1343
rect 260 1275 271 1309
rect 305 1275 316 1309
rect 260 1241 316 1275
rect 260 1207 271 1241
rect 305 1207 316 1241
rect 260 1173 316 1207
rect 260 1139 271 1173
rect 305 1139 316 1173
rect 260 1105 316 1139
rect 260 1071 271 1105
rect 305 1071 316 1105
rect 260 1037 316 1071
rect 260 1003 271 1037
rect 305 1003 316 1037
rect 260 969 316 1003
rect 260 935 271 969
rect 305 935 316 969
rect 260 865 316 935
rect 436 1853 492 1865
rect 436 1819 447 1853
rect 481 1819 492 1853
rect 436 1785 492 1819
rect 436 1751 447 1785
rect 481 1751 492 1785
rect 436 1717 492 1751
rect 436 1683 447 1717
rect 481 1683 492 1717
rect 436 1649 492 1683
rect 436 1615 447 1649
rect 481 1615 492 1649
rect 436 1581 492 1615
rect 436 1547 447 1581
rect 481 1547 492 1581
rect 436 1513 492 1547
rect 436 1479 447 1513
rect 481 1479 492 1513
rect 436 1445 492 1479
rect 436 1411 447 1445
rect 481 1411 492 1445
rect 436 1377 492 1411
rect 436 1343 447 1377
rect 481 1343 492 1377
rect 436 1309 492 1343
rect 436 1275 447 1309
rect 481 1275 492 1309
rect 436 1241 492 1275
rect 436 1207 447 1241
rect 481 1207 492 1241
rect 436 1173 492 1207
rect 436 1139 447 1173
rect 481 1139 492 1173
rect 436 1105 492 1139
rect 436 1071 447 1105
rect 481 1071 492 1105
rect 436 1037 492 1071
rect 436 1003 447 1037
rect 481 1003 492 1037
rect 436 969 492 1003
rect 436 935 447 969
rect 481 935 492 969
rect 436 865 492 935
rect 612 1853 665 1865
rect 612 1819 623 1853
rect 657 1819 665 1853
rect 612 1785 665 1819
rect 612 1751 623 1785
rect 657 1751 665 1785
rect 612 1717 665 1751
rect 612 1683 623 1717
rect 657 1683 665 1717
rect 612 1649 665 1683
rect 612 1615 623 1649
rect 657 1615 665 1649
rect 612 1581 665 1615
rect 612 1547 623 1581
rect 657 1547 665 1581
rect 612 1513 665 1547
rect 612 1479 623 1513
rect 657 1479 665 1513
rect 612 1445 665 1479
rect 612 1411 623 1445
rect 657 1411 665 1445
rect 612 1377 665 1411
rect 612 1343 623 1377
rect 657 1343 665 1377
rect 612 1309 665 1343
rect 612 1275 623 1309
rect 657 1275 665 1309
rect 612 1241 665 1275
rect 612 1207 623 1241
rect 657 1207 665 1241
rect 612 1173 665 1207
rect 612 1139 623 1173
rect 657 1139 665 1173
rect 612 1105 665 1139
rect 612 1071 623 1105
rect 657 1071 665 1105
rect 612 1037 665 1071
rect 612 1003 623 1037
rect 657 1003 665 1037
rect 612 969 665 1003
rect 612 935 623 969
rect 657 935 665 969
rect 612 865 665 935
<< mvndiffc >>
rect 115 590 149 624
rect 115 522 149 556
rect 115 454 149 488
rect 115 386 149 420
rect 115 318 149 352
rect 115 250 149 284
rect 115 182 149 216
rect 115 114 149 148
rect 291 590 325 624
rect 291 522 325 556
rect 291 454 325 488
rect 291 386 325 420
rect 291 318 325 352
rect 291 250 325 284
rect 291 182 325 216
rect 291 114 325 148
rect 467 590 501 624
rect 467 522 501 556
rect 467 454 501 488
rect 467 386 501 420
rect 467 318 501 352
rect 467 250 501 284
rect 467 182 501 216
rect 467 114 501 148
<< mvpdiffc >>
rect 95 1819 129 1853
rect 95 1751 129 1785
rect 95 1683 129 1717
rect 95 1615 129 1649
rect 95 1547 129 1581
rect 95 1479 129 1513
rect 95 1411 129 1445
rect 95 1343 129 1377
rect 95 1275 129 1309
rect 95 1207 129 1241
rect 95 1139 129 1173
rect 95 1071 129 1105
rect 95 1003 129 1037
rect 95 935 129 969
rect 271 1819 305 1853
rect 271 1751 305 1785
rect 271 1683 305 1717
rect 271 1615 305 1649
rect 271 1547 305 1581
rect 271 1479 305 1513
rect 271 1411 305 1445
rect 271 1343 305 1377
rect 271 1275 305 1309
rect 271 1207 305 1241
rect 271 1139 305 1173
rect 271 1071 305 1105
rect 271 1003 305 1037
rect 271 935 305 969
rect 447 1819 481 1853
rect 447 1751 481 1785
rect 447 1683 481 1717
rect 447 1615 481 1649
rect 447 1547 481 1581
rect 447 1479 481 1513
rect 447 1411 481 1445
rect 447 1343 481 1377
rect 447 1275 481 1309
rect 447 1207 481 1241
rect 447 1139 481 1173
rect 447 1071 481 1105
rect 447 1003 481 1037
rect 447 935 481 969
rect 623 1819 657 1853
rect 623 1751 657 1785
rect 623 1683 657 1717
rect 623 1615 657 1649
rect 623 1547 657 1581
rect 623 1479 657 1513
rect 623 1411 657 1445
rect 623 1343 657 1377
rect 623 1275 657 1309
rect 623 1207 657 1241
rect 623 1139 657 1173
rect 623 1071 657 1105
rect 623 1003 657 1037
rect 623 935 657 969
<< poly >>
rect 316 1947 612 1967
rect 316 1913 345 1947
rect 379 1913 413 1947
rect 447 1913 481 1947
rect 515 1913 549 1947
rect 583 1913 612 1947
rect 316 1891 612 1913
rect 140 1865 260 1891
rect 316 1865 436 1891
rect 492 1865 612 1891
rect 140 839 260 865
rect 316 839 436 865
rect 492 839 612 865
rect 115 803 260 839
rect 115 769 135 803
rect 169 769 203 803
rect 237 769 260 803
rect 115 728 260 769
rect 336 807 673 839
rect 336 773 551 807
rect 585 773 619 807
rect 653 773 673 807
rect 336 728 673 773
rect 160 702 280 728
rect 336 702 456 728
rect 160 76 280 102
rect 138 57 280 76
rect 138 23 158 57
rect 192 23 226 57
rect 260 23 280 57
rect 138 7 280 23
rect 336 76 456 102
rect 336 57 480 76
rect 336 23 358 57
rect 392 23 426 57
rect 460 23 480 57
rect 336 7 480 23
<< polycont >>
rect 345 1913 379 1947
rect 413 1913 447 1947
rect 481 1913 515 1947
rect 549 1913 583 1947
rect 135 769 169 803
rect 203 769 237 803
rect 551 773 585 807
rect 619 773 653 807
rect 158 23 192 57
rect 226 23 260 57
rect 358 23 392 57
rect 426 23 460 57
<< locali >>
rect 329 1913 345 1947
rect 379 1913 413 1947
rect 447 1913 481 1947
rect 515 1913 549 1947
rect 583 1913 599 1947
rect 95 1853 129 1869
rect 95 1785 129 1819
rect 95 1717 129 1751
rect 95 1649 129 1683
rect 95 1581 129 1615
rect 95 1513 129 1547
rect 95 1445 129 1479
rect 95 1377 129 1411
rect 95 1309 129 1343
rect 95 1255 129 1275
rect 271 1853 305 1869
rect 271 1785 305 1819
rect 271 1717 305 1751
rect 271 1649 305 1683
rect 271 1581 305 1615
rect 271 1513 305 1547
rect 271 1445 305 1479
rect 271 1377 305 1411
rect 271 1309 305 1343
rect 129 1221 167 1255
rect 271 1241 305 1275
rect 447 1853 481 1869
rect 447 1785 481 1819
rect 447 1717 481 1751
rect 447 1649 481 1683
rect 447 1581 481 1615
rect 447 1513 481 1547
rect 447 1445 481 1479
rect 447 1377 481 1411
rect 447 1309 481 1343
rect 447 1255 481 1275
rect 623 1853 657 1869
rect 623 1785 657 1819
rect 623 1717 657 1751
rect 623 1649 657 1683
rect 623 1581 657 1615
rect 623 1513 657 1547
rect 623 1445 657 1479
rect 623 1377 657 1411
rect 623 1309 657 1343
rect 95 1173 129 1207
rect 95 1105 129 1139
rect 95 1037 129 1071
rect 95 969 129 1003
rect 95 919 129 935
rect 443 1241 481 1255
rect 443 1221 447 1241
rect 271 1173 305 1207
rect 271 1105 305 1139
rect 271 1037 305 1067
rect 271 969 305 995
rect 271 919 305 923
rect 623 1241 657 1275
rect 447 1173 481 1207
rect 447 1105 481 1139
rect 447 1037 481 1071
rect 447 969 481 1003
rect 447 803 481 935
rect 623 1173 657 1207
rect 623 1105 657 1139
rect 623 1037 657 1067
rect 623 969 657 995
rect 623 919 657 923
rect 119 769 135 803
rect 169 769 203 803
rect 237 769 253 803
rect 447 769 501 803
rect 535 773 551 807
rect 585 773 619 807
rect 653 773 669 807
rect 115 624 149 640
rect 115 568 149 590
rect 115 496 149 522
rect 115 424 149 454
rect 115 352 149 386
rect 115 284 149 318
rect 115 216 149 250
rect 115 148 149 182
rect 115 98 149 114
rect 291 624 325 640
rect 291 556 325 590
rect 291 488 325 522
rect 291 420 325 454
rect 291 352 325 386
rect 291 284 325 318
rect 291 216 325 250
rect 291 148 325 182
rect 291 98 325 114
rect 467 624 501 769
rect 467 556 501 590
rect 467 488 501 522
rect 467 420 501 454
rect 467 352 501 386
rect 467 284 501 318
rect 467 216 501 250
rect 467 148 501 182
rect 467 98 501 114
rect 142 23 158 57
rect 192 23 226 57
rect 260 23 276 57
rect 342 23 358 57
rect 392 23 426 57
rect 460 23 476 57
<< viali >>
rect 95 1241 129 1255
rect 95 1221 129 1241
rect 167 1221 201 1255
rect 409 1221 443 1255
rect 271 1071 305 1101
rect 271 1067 305 1071
rect 271 1003 305 1029
rect 271 995 305 1003
rect 271 935 305 957
rect 271 923 305 935
rect 481 1221 515 1255
rect 623 1071 657 1101
rect 623 1067 657 1071
rect 623 1003 657 1029
rect 623 995 657 1003
rect 623 935 657 957
rect 623 923 657 935
rect 115 556 149 568
rect 115 534 149 556
rect 115 488 149 496
rect 115 462 149 488
rect 115 420 149 424
rect 115 390 149 420
<< metal1 >>
rect 83 1255 527 1261
rect 83 1221 95 1255
rect 129 1221 167 1255
rect 201 1221 409 1255
rect 443 1221 481 1255
rect 515 1221 527 1255
rect 83 1215 527 1221
rect 21 1101 731 1107
rect 21 1067 271 1101
rect 305 1067 623 1101
rect 657 1067 731 1101
rect 21 1029 731 1067
rect 21 995 271 1029
rect 305 995 623 1029
rect 657 995 731 1029
rect 21 957 731 995
rect 21 923 271 957
rect 305 923 623 957
rect 657 923 731 957
rect 21 905 731 923
rect 21 568 731 581
rect 21 534 115 568
rect 149 534 731 568
rect 21 496 731 534
rect 21 462 115 496
rect 149 462 731 496
rect 21 424 731 462
rect 21 390 115 424
rect 149 390 731 424
rect 21 379 731 390
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_0
timestamp 1663361622
transform 1 0 336 0 1 102
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_1
timestamp 1663361622
transform 1 0 160 0 1 102
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808284  sky130_fd_pr__pfet_01v8__example_55959141808284_0
timestamp 1663361622
transform -1 0 260 0 -1 1865
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808361  sky130_fd_pr__pfet_01v8__example_55959141808361_0
timestamp 1663361622
transform -1 0 612 0 -1 1865
box -1 0 297 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1663361622
transform -1 0 201 0 -1 1255
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1663361622
transform -1 0 515 0 -1 1255
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1663361622
transform 1 0 271 0 -1 1101
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1663361622
transform 1 0 623 0 -1 1101
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_2
timestamp 1663361622
transform 1 0 115 0 1 390
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1663361622
transform 0 -1 253 1 0 753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1663361622
transform 0 1 535 1 0 757
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1663361622
transform 0 -1 476 1 0 7
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1663361622
transform 0 -1 276 1 0 7
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1663361622
transform 0 1 329 1 0 1897
box 0 0 1 1
<< labels >>
flabel locali s 541 773 575 807 2 FreeSans 300 0 0 0 DRVHI_H
port 1 nsew
flabel locali s 147 769 188 803 8 FreeSans 300 0 0 0 PUEN_H
port 2 nsew
flabel metal1 s 83 1215 123 1261 3 FreeSans 300 180 0 0 PU_H_N
port 3 nsew
flabel metal1 s 21 379 63 581 7 FreeSans 300 0 0 0 VGND_IO
port 4 nsew
flabel metal1 s 689 379 731 581 7 FreeSans 300 180 0 0 VGND_IO
port 4 nsew
flabel metal1 s 21 905 58 1107 7 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 694 905 731 1107 6 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 487 1215 527 1261 3 FreeSans 300 0 0 0 PU_H_N
port 3 nsew
<< properties >>
string GDS_END 32396844
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 32393608
<< end >>
