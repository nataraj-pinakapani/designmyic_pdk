magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 74 51 75 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 74 46 75 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 7 1 12 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 12 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 7 1 11 4 VCCD
port 3 nsew power bidirectional
rlabel  s 74 7 75 11 6 VCCD
port 3 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 0 1 5 4 VCCHIB
port 4 nsew power bidirectional
rlabel  s 74 0 75 5 6 VCCHIB
port 4 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 13 1 16 4 VDDA
port 5 nsew power bidirectional
rlabel  s 74 13 75 16 6 VDDA
port 5 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 18 1 22 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 68 1 93 4 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 18 75 22 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 74 68 75 93 6 VDDIO
port 6 nsew power bidirectional
rlabel  s 0 62 1 67 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 67 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 62 1 66 4 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 74 62 75 66 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 50 1 51 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 46 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 50 75 51 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 54 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 35 1 38 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 0 46 1 55 4 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 35 75 38 6 VSSA
port 8 nsew ground bidirectional
rlabel  s 74 46 75 55 6 VSSA
port 8 nsew ground bidirectional
rlabel 
 s 1 40 25 44 6 VSSD
port 9 nsew ground bidirectional
rlabel 
 s 51 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 40 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 51 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 40 1 44 4 VSSD
port 9 nsew ground bidirectional
rlabel  s 74 40 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 75 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 75 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 75 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 75 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 75 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 75 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 75 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 75 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 40 75 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 40 75 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 74 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 74 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 40 74 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 40 74 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 44 74 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 43 74 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 42 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 74 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 74 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 41 74 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 40 74 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 74 40 74 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 41 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 41 73 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 41 73 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 40 73 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 40 73 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 41 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 41 73 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 41 73 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 40 73 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 73 40 73 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 73 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 73 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 73 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 73 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 73 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 40 73 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 40 73 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 72 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 72 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 40 72 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 40 72 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 44 72 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 43 72 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 42 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 72 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 72 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 41 72 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 40 72 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 72 40 72 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 41 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 41 71 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 41 71 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 40 71 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 40 71 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 41 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 41 71 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 41 71 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 40 71 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 71 40 71 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 71 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 71 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 71 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 71 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 71 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 40 71 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 40 71 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 70 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 70 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 40 70 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 40 70 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 44 70 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 43 70 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 42 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 70 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 70 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 41 70 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 40 70 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 70 40 70 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 41 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 41 69 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 41 69 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 40 69 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 40 69 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 41 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 41 69 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 41 69 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 40 69 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 69 40 69 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 69 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 69 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 69 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 69 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 69 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 40 69 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 40 69 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 68 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 68 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 40 68 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 40 68 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 44 68 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 43 68 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 42 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 68 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 68 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 41 68 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 40 68 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 68 40 68 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 41 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 41 67 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 41 67 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 40 67 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 40 67 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 41 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 41 67 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 41 67 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 40 67 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 67 40 67 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 67 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 67 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 67 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 67 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 67 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 40 67 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 40 67 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 66 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 66 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 40 66 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 40 66 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 44 66 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 43 66 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 42 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 66 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 66 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 41 66 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 40 66 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 66 40 66 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 41 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 41 65 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 41 65 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 40 65 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 40 65 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 44 65 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 43 65 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 42 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 41 65 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 41 65 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 41 65 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 40 65 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 65 40 65 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 41 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 41 64 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 41 64 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 40 64 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 40 64 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 41 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 41 64 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 41 64 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 40 64 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 64 40 64 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 64 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 64 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 64 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 64 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 64 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 40 64 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 40 64 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 63 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 63 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 40 63 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 40 63 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 44 63 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 43 63 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 42 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 63 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 63 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 41 63 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 40 63 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 63 40 63 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 41 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 41 62 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 41 62 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 40 62 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 40 62 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 41 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 41 62 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 41 62 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 40 62 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 62 40 62 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 62 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 62 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 62 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 62 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 62 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 40 62 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 40 62 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 61 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 61 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 40 61 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 40 61 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 44 61 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 43 61 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 42 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 61 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 61 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 41 61 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 40 61 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 61 40 61 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 41 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 41 60 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 41 60 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 40 60 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 40 60 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 41 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 41 60 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 41 60 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 40 60 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 60 40 60 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 60 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 60 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 60 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 60 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 60 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 40 60 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 40 60 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 59 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 59 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 40 59 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 40 59 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 44 59 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 43 59 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 42 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 59 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 59 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 41 59 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 40 59 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 59 40 59 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 41 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 41 58 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 41 58 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 40 58 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 40 58 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 41 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 41 58 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 41 58 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 40 58 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 58 40 58 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 58 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 58 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 58 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 58 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 58 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 40 58 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 40 58 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 57 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 57 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 40 57 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 40 57 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 44 57 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 43 57 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 42 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 57 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 57 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 41 57 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 40 57 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 57 40 57 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 41 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 41 56 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 41 56 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 40 56 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 40 56 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 41 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 41 56 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 41 56 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 40 56 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 56 40 56 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 56 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 56 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 56 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 56 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 56 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 40 56 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 40 56 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 55 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 55 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 40 55 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 40 55 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 44 55 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 43 55 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 42 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 55 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 55 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 41 55 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 40 55 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 55 40 55 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 41 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 41 54 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 41 54 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 40 54 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 40 54 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 41 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 41 54 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 41 54 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 40 54 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 54 40 54 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 54 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 54 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 41 54 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 41 54 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 41 54 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 40 54 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 40 54 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 41 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 41 53 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 41 53 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 40 53 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 53 40 53 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 53 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 53 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 53 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 53 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 53 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 40 53 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 40 53 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 52 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 52 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 40 52 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 40 52 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 44 52 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 43 52 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 42 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 52 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 52 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 41 52 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 40 52 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 52 40 52 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 41 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 41 51 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 41 51 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 40 51 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 40 51 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 44 51 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 43 51 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 42 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 41 51 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 41 51 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 41 51 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 40 51 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 51 40 51 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 41 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 41 24 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 41 24 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 40 24 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 40 24 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 41 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 41 24 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 41 24 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 40 24 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 24 40 24 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 24 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 24 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 24 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 24 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 24 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 40 24 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 40 24 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 23 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 23 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 40 23 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 40 23 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 44 23 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 43 23 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 42 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 23 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 23 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 41 23 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 40 23 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 23 40 23 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 41 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 41 22 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 41 22 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 40 22 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 40 22 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 41 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 41 22 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 41 22 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 40 22 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 22 40 22 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 22 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 22 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 22 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 22 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 22 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 40 22 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 40 22 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 21 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 21 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 40 21 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 40 21 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 44 21 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 43 21 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 42 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 21 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 21 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 41 21 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 40 21 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 21 40 21 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 41 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 41 20 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 41 20 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 40 20 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 40 20 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 41 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 41 20 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 41 20 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 40 20 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 20 40 20 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 20 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 20 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 20 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 20 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 20 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 40 20 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 40 20 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 19 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 19 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 40 19 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 40 19 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 44 19 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 43 19 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 42 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 19 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 19 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 41 19 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 40 19 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 19 40 19 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 41 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 41 18 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 41 18 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 40 18 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 40 18 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 41 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 41 18 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 41 18 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 40 18 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 18 40 18 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 18 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 18 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 18 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 18 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 18 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 40 18 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 40 18 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 17 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 17 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 40 17 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 40 17 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 44 17 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 43 17 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 42 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 17 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 17 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 41 17 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 40 17 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 17 40 17 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 41 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 41 16 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 41 16 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 40 16 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 40 16 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 41 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 41 16 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 41 16 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 40 16 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 16 40 16 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 16 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 16 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 16 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 16 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 16 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 40 16 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 40 16 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 15 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 15 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 40 15 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 40 15 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 44 15 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 43 15 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 42 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 15 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 15 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 41 15 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 40 15 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 15 40 15 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 41 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 41 14 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 41 14 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 40 14 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 40 14 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 41 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 41 14 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 41 14 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 40 14 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 14 40 14 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 14 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 14 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 14 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 14 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 14 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 40 14 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 40 14 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 13 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 13 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 40 13 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 40 13 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 44 13 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 43 13 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 42 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 13 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 13 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 41 13 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 40 13 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 13 40 13 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 41 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 41 12 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 41 12 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 40 12 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 40 12 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 41 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 41 12 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 41 12 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 40 12 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 12 40 12 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 12 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 12 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 12 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 12 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 12 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 40 12 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 40 12 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 11 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 11 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 40 11 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 40 11 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 44 11 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 43 11 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 42 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 11 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 11 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 41 11 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 40 11 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 11 40 11 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 41 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 41 10 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 41 10 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 40 10 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 40 10 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 41 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 41 10 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 41 10 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 40 10 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 10 40 10 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 10 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 10 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 10 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 10 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 10 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 40 10 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 40 10 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 9 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 9 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 40 9 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 40 9 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 44 9 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 43 9 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 42 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 9 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 9 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 41 9 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 40 9 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 9 40 9 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 41 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 41 8 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 41 8 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 40 8 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 40 8 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 41 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 41 8 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 41 8 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 40 8 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 8 40 8 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 8 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 8 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 8 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 8 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 8 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 40 8 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 40 8 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 7 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 7 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 40 7 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 40 7 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 44 7 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 43 7 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 42 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 7 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 7 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 41 7 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 40 7 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 7 40 7 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 41 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 41 6 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 41 6 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 40 6 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 40 6 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 41 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 41 6 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 41 6 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 40 6 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 6 40 6 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 6 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 6 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 6 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 6 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 6 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 40 6 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 40 6 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 5 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 5 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 40 5 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 40 5 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 44 5 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 43 5 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 42 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 5 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 5 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 41 5 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 40 5 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 5 40 5 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 41 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 41 4 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 41 4 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 40 4 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 40 4 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 41 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 41 4 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 41 4 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 40 4 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 4 40 4 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 4 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 4 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 4 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 4 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 4 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 40 4 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 40 4 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 3 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 3 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 40 3 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 40 3 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 44 3 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 43 3 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 42 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 3 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 3 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 41 3 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 40 3 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 3 40 3 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 41 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 41 2 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 41 2 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 40 2 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 40 2 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 41 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 41 2 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 41 2 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 40 2 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 2 40 2 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 2 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 2 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 2 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 2 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 2 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 40 2 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 40 2 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 1 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 1 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 1 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 1 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 1 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 1 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 40 1 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 40 1 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 1 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 44 1 44 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 1 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 43 1 43 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 42 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 1 42 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 1 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 41 1 41 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 40 1 40 6 VSSD
port 9 nsew ground bidirectional
rlabel nfet_brown s 1 40 1 40 6 VSSD
port 9 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 24 1 28 4 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 174 75 198 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 74 24 75 28 6 VSSIO
port 10 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 56 1 61 4 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 74 56 75 61 6 VSSIO_Q
port 11 nsew ground bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
rlabel  s 0 30 1 33 4 VSWITCH
port 12 nsew power bidirectional
rlabel  s 74 30 75 33 6 VSWITCH
port 12 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 75 198
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
