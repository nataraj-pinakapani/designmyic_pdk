magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 11 21 905 203
rect 25 -17 59 21
<< scnmos >>
rect 90 47 120 177
rect 176 47 206 177
rect 262 47 292 177
rect 348 47 378 177
rect 538 47 568 177
rect 624 47 654 177
rect 710 47 740 177
rect 796 47 826 177
<< scpmoshvt >>
rect 90 297 120 497
rect 176 297 206 497
rect 262 297 292 497
rect 348 297 378 497
rect 538 297 568 497
rect 624 297 654 497
rect 710 297 740 497
rect 796 297 826 497
<< ndiff >>
rect 37 135 90 177
rect 37 101 45 135
rect 79 101 90 135
rect 37 47 90 101
rect 120 169 176 177
rect 120 135 131 169
rect 165 135 176 169
rect 120 101 176 135
rect 120 67 131 101
rect 165 67 176 101
rect 120 47 176 67
rect 206 93 262 177
rect 206 59 217 93
rect 251 59 262 93
rect 206 47 262 59
rect 292 131 348 177
rect 292 97 303 131
rect 337 97 348 131
rect 292 47 348 97
rect 378 93 431 177
rect 378 59 389 93
rect 423 59 431 93
rect 378 47 431 59
rect 485 93 538 177
rect 485 59 493 93
rect 527 59 538 93
rect 485 47 538 59
rect 568 168 624 177
rect 568 134 579 168
rect 613 134 624 168
rect 568 47 624 134
rect 654 124 710 177
rect 654 90 665 124
rect 699 90 710 124
rect 654 47 710 90
rect 740 89 796 177
rect 740 55 751 89
rect 785 55 796 89
rect 740 47 796 55
rect 826 127 879 177
rect 826 93 837 127
rect 871 93 879 127
rect 826 47 879 93
<< pdiff >>
rect 37 475 90 497
rect 37 441 45 475
rect 79 441 90 475
rect 37 407 90 441
rect 37 373 45 407
rect 79 373 90 407
rect 37 297 90 373
rect 120 415 176 497
rect 120 381 131 415
rect 165 381 176 415
rect 120 347 176 381
rect 120 313 131 347
rect 165 313 176 347
rect 120 297 176 313
rect 206 475 262 497
rect 206 441 217 475
rect 251 441 262 475
rect 206 407 262 441
rect 206 373 217 407
rect 251 373 262 407
rect 206 297 262 373
rect 292 415 348 497
rect 292 381 303 415
rect 337 381 348 415
rect 292 347 348 381
rect 292 313 303 347
rect 337 313 348 347
rect 292 297 348 313
rect 378 485 431 497
rect 378 451 389 485
rect 423 451 431 485
rect 378 417 431 451
rect 378 383 389 417
rect 423 383 431 417
rect 378 297 431 383
rect 485 485 538 497
rect 485 451 493 485
rect 527 451 538 485
rect 485 417 538 451
rect 485 383 493 417
rect 527 383 538 417
rect 485 297 538 383
rect 568 477 624 497
rect 568 443 579 477
rect 613 443 624 477
rect 568 409 624 443
rect 568 375 579 409
rect 613 375 624 409
rect 568 341 624 375
rect 568 307 579 341
rect 613 307 624 341
rect 568 297 624 307
rect 654 485 710 497
rect 654 451 665 485
rect 699 451 710 485
rect 654 417 710 451
rect 654 383 665 417
rect 699 383 710 417
rect 654 297 710 383
rect 740 477 796 497
rect 740 443 751 477
rect 785 443 796 477
rect 740 409 796 443
rect 740 375 751 409
rect 785 375 796 409
rect 740 341 796 375
rect 740 307 751 341
rect 785 307 796 341
rect 740 297 796 307
rect 826 485 879 497
rect 826 451 837 485
rect 871 451 879 485
rect 826 417 879 451
rect 826 383 837 417
rect 871 383 879 417
rect 826 297 879 383
<< ndiffc >>
rect 45 101 79 135
rect 131 135 165 169
rect 131 67 165 101
rect 217 59 251 93
rect 303 97 337 131
rect 389 59 423 93
rect 493 59 527 93
rect 579 134 613 168
rect 665 90 699 124
rect 751 55 785 89
rect 837 93 871 127
<< pdiffc >>
rect 45 441 79 475
rect 45 373 79 407
rect 131 381 165 415
rect 131 313 165 347
rect 217 441 251 475
rect 217 373 251 407
rect 303 381 337 415
rect 303 313 337 347
rect 389 451 423 485
rect 389 383 423 417
rect 493 451 527 485
rect 493 383 527 417
rect 579 443 613 477
rect 579 375 613 409
rect 579 307 613 341
rect 665 451 699 485
rect 665 383 699 417
rect 751 443 785 477
rect 751 375 785 409
rect 751 307 785 341
rect 837 451 871 485
rect 837 383 871 417
<< poly >>
rect 90 497 120 523
rect 176 497 206 523
rect 262 497 292 523
rect 348 497 378 523
rect 538 497 568 523
rect 624 497 654 523
rect 710 497 740 523
rect 796 497 826 523
rect 90 265 120 297
rect 176 265 206 297
rect 36 249 206 265
rect 36 215 46 249
rect 80 215 206 249
rect 36 199 206 215
rect 90 177 120 199
rect 176 177 206 199
rect 262 265 292 297
rect 348 265 378 297
rect 538 265 568 297
rect 624 265 654 297
rect 262 249 378 265
rect 262 215 303 249
rect 337 215 378 249
rect 262 199 378 215
rect 484 249 654 265
rect 484 215 494 249
rect 528 215 562 249
rect 596 215 654 249
rect 484 199 654 215
rect 262 177 292 199
rect 348 177 378 199
rect 538 177 568 199
rect 624 177 654 199
rect 710 265 740 297
rect 796 265 826 297
rect 710 249 880 265
rect 710 215 768 249
rect 802 215 836 249
rect 870 215 880 249
rect 710 199 880 215
rect 710 177 740 199
rect 796 177 826 199
rect 90 21 120 47
rect 176 21 206 47
rect 262 21 292 47
rect 348 21 378 47
rect 538 21 568 47
rect 624 21 654 47
rect 710 21 740 47
rect 796 21 826 47
<< polycont >>
rect 46 215 80 249
rect 303 215 337 249
rect 494 215 528 249
rect 562 215 596 249
rect 768 215 802 249
rect 836 215 870 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 29 485 443 491
rect 29 475 389 485
rect 29 441 45 475
rect 79 457 217 475
rect 79 441 81 457
rect 29 407 81 441
rect 215 441 217 457
rect 251 451 389 475
rect 423 451 443 485
rect 251 441 253 451
rect 29 373 45 407
rect 79 373 81 407
rect 29 357 81 373
rect 115 415 181 421
rect 115 381 131 415
rect 165 381 181 415
rect 115 357 181 381
rect 215 407 253 441
rect 387 417 443 451
rect 215 373 217 407
rect 251 373 253 407
rect 215 357 253 373
rect 287 381 303 415
rect 337 381 353 415
rect 115 347 171 357
rect 20 249 81 323
rect 20 215 46 249
rect 80 215 81 249
rect 20 199 81 215
rect 115 313 131 347
rect 165 313 171 347
rect 287 347 353 381
rect 387 383 389 417
rect 423 383 443 417
rect 387 367 443 383
rect 487 485 533 527
rect 487 451 493 485
rect 527 451 533 485
rect 487 417 533 451
rect 487 383 493 417
rect 527 383 533 417
rect 487 367 533 383
rect 569 477 623 493
rect 569 443 579 477
rect 613 443 623 477
rect 569 409 623 443
rect 569 375 579 409
rect 613 375 623 409
rect 115 171 171 313
rect 207 257 251 323
rect 287 313 303 347
rect 337 331 353 347
rect 569 341 623 375
rect 659 485 705 527
rect 659 451 665 485
rect 699 451 705 485
rect 659 417 705 451
rect 659 383 665 417
rect 699 383 705 417
rect 659 367 705 383
rect 741 477 795 493
rect 741 443 751 477
rect 785 443 795 477
rect 741 409 795 443
rect 741 375 751 409
rect 785 375 795 409
rect 569 331 579 341
rect 337 313 579 331
rect 287 307 579 313
rect 613 331 623 341
rect 741 341 795 375
rect 831 485 877 527
rect 831 451 837 485
rect 871 451 877 485
rect 831 417 877 451
rect 831 383 837 417
rect 871 383 877 417
rect 831 367 877 383
rect 741 331 751 341
rect 613 307 751 331
rect 785 307 795 341
rect 287 291 795 307
rect 835 257 900 331
rect 207 249 357 257
rect 207 215 303 249
rect 337 215 357 249
rect 207 207 357 215
rect 474 249 616 257
rect 474 215 494 249
rect 528 215 562 249
rect 596 215 616 249
rect 474 207 616 215
rect 748 249 900 257
rect 748 215 768 249
rect 802 215 836 249
rect 870 215 900 249
rect 748 207 900 215
rect 115 169 629 171
rect 29 135 79 163
rect 29 101 45 135
rect 29 17 79 101
rect 115 135 131 169
rect 165 168 629 169
rect 165 135 579 168
rect 115 134 579 135
rect 613 134 629 168
rect 115 131 629 134
rect 115 101 167 131
rect 115 67 131 101
rect 165 67 167 101
rect 301 97 303 131
rect 337 97 339 131
rect 115 51 167 67
rect 201 93 267 95
rect 201 59 217 93
rect 251 59 267 93
rect 201 17 267 59
rect 301 57 339 97
rect 665 127 887 171
rect 665 124 699 127
rect 373 93 439 95
rect 373 59 389 93
rect 423 59 439 93
rect 373 17 439 59
rect 477 93 665 95
rect 477 59 493 93
rect 527 90 665 93
rect 871 93 887 127
rect 527 59 699 90
rect 477 53 699 59
rect 735 89 801 91
rect 735 55 751 89
rect 785 55 801 89
rect 735 17 801 55
rect 837 53 887 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 765 221 799 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 25 221 59 255 0 FreeSans 200 0 0 0 C1
port 4 nsew signal input
flabel locali s 25 289 59 323 0 FreeSans 200 0 0 0 C1
port 4 nsew signal input
flabel locali s 301 221 335 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 117 289 151 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 117 357 151 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 117 221 151 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 117 153 151 187 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 117 85 151 119 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 301 85 335 119 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 857 289 891 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 209 221 243 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 209 289 243 323 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel metal1 s 25 527 59 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 25 -17 59 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 25 527 59 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 25 -17 59 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a211oi_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 3613130
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3604188
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 23.000 13.600 
<< end >>
