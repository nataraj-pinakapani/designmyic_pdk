/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__rf_nfet_01v8_lvt_cM04W5p00L0p18.spice