* SKY130 Spice File.
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_01v8__fs.pm3.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_01v8_lvt__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_03v3_nvt__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_05v0_nvt__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__esd_nfet_01v8__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8_lvt__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8_hvt__fs.pm3.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__esd_pfet_g5v0d10v5__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_g5v0d10v5__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_g5v0d16v0__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_g5v0d10v5__fs.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_g5v0d16v0__fs_discrete.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__esd_nfet_g5v0d10v5__fs.corner.spice"
.include "fs/nonfet.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_20v0__fs_discrete.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_20v0__fs_discrete.corner.spice"
.include "../../../libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_20v0_nvt__fs_discrete.corner.spice"
.include "../all.spice"
.include "fs/rf.spice"
