magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 0 2336 4043 3048
rect 0 1799 3192 2336
<< pwell >>
rect 4338 224 5304 239
rect 10 -828 5742 224
rect 41 -938 5717 -828
<< mvnmos >>
rect 89 -802 249 198
rect 305 -802 465 198
rect 521 -802 681 198
rect 737 -802 897 198
rect 953 -802 1113 198
rect 1169 -802 1329 198
rect 1385 -802 1545 198
rect 1601 -802 1761 198
rect 1817 -802 1977 198
rect 2033 -802 2193 198
rect 2249 -802 2409 198
rect 2465 -802 2625 198
rect 2681 -802 2841 198
rect 2897 -802 3057 198
rect 3113 -802 3273 198
rect 3439 -802 3599 198
rect 3765 -802 3925 198
rect 4091 -802 4251 198
rect 4417 13 4577 213
rect 4633 13 4793 213
rect 4849 13 5009 213
rect 5065 13 5225 213
rect 4417 -802 4617 -202
rect 4673 -802 4773 -202
rect 4829 -802 4929 -202
rect 4985 -802 5085 -202
rect 5141 -802 5241 -202
rect 5407 -802 5507 198
rect 5563 -802 5663 198
<< mvpmos >>
rect 119 1865 219 2865
rect 275 1865 375 2865
rect 541 1865 701 2865
rect 757 1865 917 2865
rect 973 1865 1073 2865
rect 1129 1865 1229 2865
rect 1445 1865 1605 2865
rect 1661 1865 1761 2865
rect 1817 1865 1917 2865
rect 1973 1865 2073 2865
rect 2129 1865 2229 2865
rect 2285 1865 2385 2865
rect 2551 1865 2651 2465
rect 2817 1865 2917 2865
rect 2973 1865 3073 2865
<< mvndiff >>
rect 4364 201 4417 213
rect 36 128 89 198
rect 36 94 44 128
rect 78 94 89 128
rect 36 60 89 94
rect 36 26 44 60
rect 78 26 89 60
rect 36 -8 89 26
rect 36 -42 44 -8
rect 78 -42 89 -8
rect 36 -76 89 -42
rect 36 -110 44 -76
rect 78 -110 89 -76
rect 36 -144 89 -110
rect 36 -178 44 -144
rect 78 -178 89 -144
rect 36 -212 89 -178
rect 36 -246 44 -212
rect 78 -246 89 -212
rect 36 -280 89 -246
rect 36 -314 44 -280
rect 78 -314 89 -280
rect 36 -348 89 -314
rect 36 -382 44 -348
rect 78 -382 89 -348
rect 36 -416 89 -382
rect 36 -450 44 -416
rect 78 -450 89 -416
rect 36 -484 89 -450
rect 36 -518 44 -484
rect 78 -518 89 -484
rect 36 -552 89 -518
rect 36 -586 44 -552
rect 78 -586 89 -552
rect 36 -620 89 -586
rect 36 -654 44 -620
rect 78 -654 89 -620
rect 36 -688 89 -654
rect 36 -722 44 -688
rect 78 -722 89 -688
rect 36 -756 89 -722
rect 36 -790 44 -756
rect 78 -790 89 -756
rect 36 -802 89 -790
rect 249 128 305 198
rect 249 94 260 128
rect 294 94 305 128
rect 249 60 305 94
rect 249 26 260 60
rect 294 26 305 60
rect 249 -8 305 26
rect 249 -42 260 -8
rect 294 -42 305 -8
rect 249 -76 305 -42
rect 249 -110 260 -76
rect 294 -110 305 -76
rect 249 -144 305 -110
rect 249 -178 260 -144
rect 294 -178 305 -144
rect 249 -212 305 -178
rect 249 -246 260 -212
rect 294 -246 305 -212
rect 249 -280 305 -246
rect 249 -314 260 -280
rect 294 -314 305 -280
rect 249 -348 305 -314
rect 249 -382 260 -348
rect 294 -382 305 -348
rect 249 -416 305 -382
rect 249 -450 260 -416
rect 294 -450 305 -416
rect 249 -484 305 -450
rect 249 -518 260 -484
rect 294 -518 305 -484
rect 249 -552 305 -518
rect 249 -586 260 -552
rect 294 -586 305 -552
rect 249 -620 305 -586
rect 249 -654 260 -620
rect 294 -654 305 -620
rect 249 -688 305 -654
rect 249 -722 260 -688
rect 294 -722 305 -688
rect 249 -756 305 -722
rect 249 -790 260 -756
rect 294 -790 305 -756
rect 249 -802 305 -790
rect 465 128 521 198
rect 465 94 476 128
rect 510 94 521 128
rect 465 60 521 94
rect 465 26 476 60
rect 510 26 521 60
rect 465 -8 521 26
rect 465 -42 476 -8
rect 510 -42 521 -8
rect 465 -76 521 -42
rect 465 -110 476 -76
rect 510 -110 521 -76
rect 465 -144 521 -110
rect 465 -178 476 -144
rect 510 -178 521 -144
rect 465 -212 521 -178
rect 465 -246 476 -212
rect 510 -246 521 -212
rect 465 -280 521 -246
rect 465 -314 476 -280
rect 510 -314 521 -280
rect 465 -348 521 -314
rect 465 -382 476 -348
rect 510 -382 521 -348
rect 465 -416 521 -382
rect 465 -450 476 -416
rect 510 -450 521 -416
rect 465 -484 521 -450
rect 465 -518 476 -484
rect 510 -518 521 -484
rect 465 -552 521 -518
rect 465 -586 476 -552
rect 510 -586 521 -552
rect 465 -620 521 -586
rect 465 -654 476 -620
rect 510 -654 521 -620
rect 465 -688 521 -654
rect 465 -722 476 -688
rect 510 -722 521 -688
rect 465 -756 521 -722
rect 465 -790 476 -756
rect 510 -790 521 -756
rect 465 -802 521 -790
rect 681 128 737 198
rect 681 94 692 128
rect 726 94 737 128
rect 681 60 737 94
rect 681 26 692 60
rect 726 26 737 60
rect 681 -8 737 26
rect 681 -42 692 -8
rect 726 -42 737 -8
rect 681 -76 737 -42
rect 681 -110 692 -76
rect 726 -110 737 -76
rect 681 -144 737 -110
rect 681 -178 692 -144
rect 726 -178 737 -144
rect 681 -212 737 -178
rect 681 -246 692 -212
rect 726 -246 737 -212
rect 681 -280 737 -246
rect 681 -314 692 -280
rect 726 -314 737 -280
rect 681 -348 737 -314
rect 681 -382 692 -348
rect 726 -382 737 -348
rect 681 -416 737 -382
rect 681 -450 692 -416
rect 726 -450 737 -416
rect 681 -484 737 -450
rect 681 -518 692 -484
rect 726 -518 737 -484
rect 681 -552 737 -518
rect 681 -586 692 -552
rect 726 -586 737 -552
rect 681 -620 737 -586
rect 681 -654 692 -620
rect 726 -654 737 -620
rect 681 -688 737 -654
rect 681 -722 692 -688
rect 726 -722 737 -688
rect 681 -756 737 -722
rect 681 -790 692 -756
rect 726 -790 737 -756
rect 681 -802 737 -790
rect 897 128 953 198
rect 897 94 908 128
rect 942 94 953 128
rect 897 60 953 94
rect 897 26 908 60
rect 942 26 953 60
rect 897 -8 953 26
rect 897 -42 908 -8
rect 942 -42 953 -8
rect 897 -76 953 -42
rect 897 -110 908 -76
rect 942 -110 953 -76
rect 897 -144 953 -110
rect 897 -178 908 -144
rect 942 -178 953 -144
rect 897 -212 953 -178
rect 897 -246 908 -212
rect 942 -246 953 -212
rect 897 -280 953 -246
rect 897 -314 908 -280
rect 942 -314 953 -280
rect 897 -348 953 -314
rect 897 -382 908 -348
rect 942 -382 953 -348
rect 897 -416 953 -382
rect 897 -450 908 -416
rect 942 -450 953 -416
rect 897 -484 953 -450
rect 897 -518 908 -484
rect 942 -518 953 -484
rect 897 -552 953 -518
rect 897 -586 908 -552
rect 942 -586 953 -552
rect 897 -620 953 -586
rect 897 -654 908 -620
rect 942 -654 953 -620
rect 897 -688 953 -654
rect 897 -722 908 -688
rect 942 -722 953 -688
rect 897 -756 953 -722
rect 897 -790 908 -756
rect 942 -790 953 -756
rect 897 -802 953 -790
rect 1113 128 1169 198
rect 1113 94 1124 128
rect 1158 94 1169 128
rect 1113 60 1169 94
rect 1113 26 1124 60
rect 1158 26 1169 60
rect 1113 -8 1169 26
rect 1113 -42 1124 -8
rect 1158 -42 1169 -8
rect 1113 -76 1169 -42
rect 1113 -110 1124 -76
rect 1158 -110 1169 -76
rect 1113 -144 1169 -110
rect 1113 -178 1124 -144
rect 1158 -178 1169 -144
rect 1113 -212 1169 -178
rect 1113 -246 1124 -212
rect 1158 -246 1169 -212
rect 1113 -280 1169 -246
rect 1113 -314 1124 -280
rect 1158 -314 1169 -280
rect 1113 -348 1169 -314
rect 1113 -382 1124 -348
rect 1158 -382 1169 -348
rect 1113 -416 1169 -382
rect 1113 -450 1124 -416
rect 1158 -450 1169 -416
rect 1113 -484 1169 -450
rect 1113 -518 1124 -484
rect 1158 -518 1169 -484
rect 1113 -552 1169 -518
rect 1113 -586 1124 -552
rect 1158 -586 1169 -552
rect 1113 -620 1169 -586
rect 1113 -654 1124 -620
rect 1158 -654 1169 -620
rect 1113 -688 1169 -654
rect 1113 -722 1124 -688
rect 1158 -722 1169 -688
rect 1113 -756 1169 -722
rect 1113 -790 1124 -756
rect 1158 -790 1169 -756
rect 1113 -802 1169 -790
rect 1329 128 1385 198
rect 1329 94 1340 128
rect 1374 94 1385 128
rect 1329 60 1385 94
rect 1329 26 1340 60
rect 1374 26 1385 60
rect 1329 -8 1385 26
rect 1329 -42 1340 -8
rect 1374 -42 1385 -8
rect 1329 -76 1385 -42
rect 1329 -110 1340 -76
rect 1374 -110 1385 -76
rect 1329 -144 1385 -110
rect 1329 -178 1340 -144
rect 1374 -178 1385 -144
rect 1329 -212 1385 -178
rect 1329 -246 1340 -212
rect 1374 -246 1385 -212
rect 1329 -280 1385 -246
rect 1329 -314 1340 -280
rect 1374 -314 1385 -280
rect 1329 -348 1385 -314
rect 1329 -382 1340 -348
rect 1374 -382 1385 -348
rect 1329 -416 1385 -382
rect 1329 -450 1340 -416
rect 1374 -450 1385 -416
rect 1329 -484 1385 -450
rect 1329 -518 1340 -484
rect 1374 -518 1385 -484
rect 1329 -552 1385 -518
rect 1329 -586 1340 -552
rect 1374 -586 1385 -552
rect 1329 -620 1385 -586
rect 1329 -654 1340 -620
rect 1374 -654 1385 -620
rect 1329 -688 1385 -654
rect 1329 -722 1340 -688
rect 1374 -722 1385 -688
rect 1329 -756 1385 -722
rect 1329 -790 1340 -756
rect 1374 -790 1385 -756
rect 1329 -802 1385 -790
rect 1545 128 1601 198
rect 1545 94 1556 128
rect 1590 94 1601 128
rect 1545 60 1601 94
rect 1545 26 1556 60
rect 1590 26 1601 60
rect 1545 -8 1601 26
rect 1545 -42 1556 -8
rect 1590 -42 1601 -8
rect 1545 -76 1601 -42
rect 1545 -110 1556 -76
rect 1590 -110 1601 -76
rect 1545 -144 1601 -110
rect 1545 -178 1556 -144
rect 1590 -178 1601 -144
rect 1545 -212 1601 -178
rect 1545 -246 1556 -212
rect 1590 -246 1601 -212
rect 1545 -280 1601 -246
rect 1545 -314 1556 -280
rect 1590 -314 1601 -280
rect 1545 -348 1601 -314
rect 1545 -382 1556 -348
rect 1590 -382 1601 -348
rect 1545 -416 1601 -382
rect 1545 -450 1556 -416
rect 1590 -450 1601 -416
rect 1545 -484 1601 -450
rect 1545 -518 1556 -484
rect 1590 -518 1601 -484
rect 1545 -552 1601 -518
rect 1545 -586 1556 -552
rect 1590 -586 1601 -552
rect 1545 -620 1601 -586
rect 1545 -654 1556 -620
rect 1590 -654 1601 -620
rect 1545 -688 1601 -654
rect 1545 -722 1556 -688
rect 1590 -722 1601 -688
rect 1545 -756 1601 -722
rect 1545 -790 1556 -756
rect 1590 -790 1601 -756
rect 1545 -802 1601 -790
rect 1761 128 1817 198
rect 1761 94 1772 128
rect 1806 94 1817 128
rect 1761 60 1817 94
rect 1761 26 1772 60
rect 1806 26 1817 60
rect 1761 -8 1817 26
rect 1761 -42 1772 -8
rect 1806 -42 1817 -8
rect 1761 -76 1817 -42
rect 1761 -110 1772 -76
rect 1806 -110 1817 -76
rect 1761 -144 1817 -110
rect 1761 -178 1772 -144
rect 1806 -178 1817 -144
rect 1761 -212 1817 -178
rect 1761 -246 1772 -212
rect 1806 -246 1817 -212
rect 1761 -280 1817 -246
rect 1761 -314 1772 -280
rect 1806 -314 1817 -280
rect 1761 -348 1817 -314
rect 1761 -382 1772 -348
rect 1806 -382 1817 -348
rect 1761 -416 1817 -382
rect 1761 -450 1772 -416
rect 1806 -450 1817 -416
rect 1761 -484 1817 -450
rect 1761 -518 1772 -484
rect 1806 -518 1817 -484
rect 1761 -552 1817 -518
rect 1761 -586 1772 -552
rect 1806 -586 1817 -552
rect 1761 -620 1817 -586
rect 1761 -654 1772 -620
rect 1806 -654 1817 -620
rect 1761 -688 1817 -654
rect 1761 -722 1772 -688
rect 1806 -722 1817 -688
rect 1761 -756 1817 -722
rect 1761 -790 1772 -756
rect 1806 -790 1817 -756
rect 1761 -802 1817 -790
rect 1977 128 2033 198
rect 1977 94 1988 128
rect 2022 94 2033 128
rect 1977 60 2033 94
rect 1977 26 1988 60
rect 2022 26 2033 60
rect 1977 -8 2033 26
rect 1977 -42 1988 -8
rect 2022 -42 2033 -8
rect 1977 -76 2033 -42
rect 1977 -110 1988 -76
rect 2022 -110 2033 -76
rect 1977 -144 2033 -110
rect 1977 -178 1988 -144
rect 2022 -178 2033 -144
rect 1977 -212 2033 -178
rect 1977 -246 1988 -212
rect 2022 -246 2033 -212
rect 1977 -280 2033 -246
rect 1977 -314 1988 -280
rect 2022 -314 2033 -280
rect 1977 -348 2033 -314
rect 1977 -382 1988 -348
rect 2022 -382 2033 -348
rect 1977 -416 2033 -382
rect 1977 -450 1988 -416
rect 2022 -450 2033 -416
rect 1977 -484 2033 -450
rect 1977 -518 1988 -484
rect 2022 -518 2033 -484
rect 1977 -552 2033 -518
rect 1977 -586 1988 -552
rect 2022 -586 2033 -552
rect 1977 -620 2033 -586
rect 1977 -654 1988 -620
rect 2022 -654 2033 -620
rect 1977 -688 2033 -654
rect 1977 -722 1988 -688
rect 2022 -722 2033 -688
rect 1977 -756 2033 -722
rect 1977 -790 1988 -756
rect 2022 -790 2033 -756
rect 1977 -802 2033 -790
rect 2193 128 2249 198
rect 2193 94 2204 128
rect 2238 94 2249 128
rect 2193 60 2249 94
rect 2193 26 2204 60
rect 2238 26 2249 60
rect 2193 -8 2249 26
rect 2193 -42 2204 -8
rect 2238 -42 2249 -8
rect 2193 -76 2249 -42
rect 2193 -110 2204 -76
rect 2238 -110 2249 -76
rect 2193 -144 2249 -110
rect 2193 -178 2204 -144
rect 2238 -178 2249 -144
rect 2193 -212 2249 -178
rect 2193 -246 2204 -212
rect 2238 -246 2249 -212
rect 2193 -280 2249 -246
rect 2193 -314 2204 -280
rect 2238 -314 2249 -280
rect 2193 -348 2249 -314
rect 2193 -382 2204 -348
rect 2238 -382 2249 -348
rect 2193 -416 2249 -382
rect 2193 -450 2204 -416
rect 2238 -450 2249 -416
rect 2193 -484 2249 -450
rect 2193 -518 2204 -484
rect 2238 -518 2249 -484
rect 2193 -552 2249 -518
rect 2193 -586 2204 -552
rect 2238 -586 2249 -552
rect 2193 -620 2249 -586
rect 2193 -654 2204 -620
rect 2238 -654 2249 -620
rect 2193 -688 2249 -654
rect 2193 -722 2204 -688
rect 2238 -722 2249 -688
rect 2193 -756 2249 -722
rect 2193 -790 2204 -756
rect 2238 -790 2249 -756
rect 2193 -802 2249 -790
rect 2409 128 2465 198
rect 2409 94 2420 128
rect 2454 94 2465 128
rect 2409 60 2465 94
rect 2409 26 2420 60
rect 2454 26 2465 60
rect 2409 -8 2465 26
rect 2409 -42 2420 -8
rect 2454 -42 2465 -8
rect 2409 -76 2465 -42
rect 2409 -110 2420 -76
rect 2454 -110 2465 -76
rect 2409 -144 2465 -110
rect 2409 -178 2420 -144
rect 2454 -178 2465 -144
rect 2409 -212 2465 -178
rect 2409 -246 2420 -212
rect 2454 -246 2465 -212
rect 2409 -280 2465 -246
rect 2409 -314 2420 -280
rect 2454 -314 2465 -280
rect 2409 -348 2465 -314
rect 2409 -382 2420 -348
rect 2454 -382 2465 -348
rect 2409 -416 2465 -382
rect 2409 -450 2420 -416
rect 2454 -450 2465 -416
rect 2409 -484 2465 -450
rect 2409 -518 2420 -484
rect 2454 -518 2465 -484
rect 2409 -552 2465 -518
rect 2409 -586 2420 -552
rect 2454 -586 2465 -552
rect 2409 -620 2465 -586
rect 2409 -654 2420 -620
rect 2454 -654 2465 -620
rect 2409 -688 2465 -654
rect 2409 -722 2420 -688
rect 2454 -722 2465 -688
rect 2409 -756 2465 -722
rect 2409 -790 2420 -756
rect 2454 -790 2465 -756
rect 2409 -802 2465 -790
rect 2625 128 2681 198
rect 2625 94 2636 128
rect 2670 94 2681 128
rect 2625 60 2681 94
rect 2625 26 2636 60
rect 2670 26 2681 60
rect 2625 -8 2681 26
rect 2625 -42 2636 -8
rect 2670 -42 2681 -8
rect 2625 -76 2681 -42
rect 2625 -110 2636 -76
rect 2670 -110 2681 -76
rect 2625 -144 2681 -110
rect 2625 -178 2636 -144
rect 2670 -178 2681 -144
rect 2625 -212 2681 -178
rect 2625 -246 2636 -212
rect 2670 -246 2681 -212
rect 2625 -280 2681 -246
rect 2625 -314 2636 -280
rect 2670 -314 2681 -280
rect 2625 -348 2681 -314
rect 2625 -382 2636 -348
rect 2670 -382 2681 -348
rect 2625 -416 2681 -382
rect 2625 -450 2636 -416
rect 2670 -450 2681 -416
rect 2625 -484 2681 -450
rect 2625 -518 2636 -484
rect 2670 -518 2681 -484
rect 2625 -552 2681 -518
rect 2625 -586 2636 -552
rect 2670 -586 2681 -552
rect 2625 -620 2681 -586
rect 2625 -654 2636 -620
rect 2670 -654 2681 -620
rect 2625 -688 2681 -654
rect 2625 -722 2636 -688
rect 2670 -722 2681 -688
rect 2625 -756 2681 -722
rect 2625 -790 2636 -756
rect 2670 -790 2681 -756
rect 2625 -802 2681 -790
rect 2841 128 2897 198
rect 2841 94 2852 128
rect 2886 94 2897 128
rect 2841 60 2897 94
rect 2841 26 2852 60
rect 2886 26 2897 60
rect 2841 -8 2897 26
rect 2841 -42 2852 -8
rect 2886 -42 2897 -8
rect 2841 -76 2897 -42
rect 2841 -110 2852 -76
rect 2886 -110 2897 -76
rect 2841 -144 2897 -110
rect 2841 -178 2852 -144
rect 2886 -178 2897 -144
rect 2841 -212 2897 -178
rect 2841 -246 2852 -212
rect 2886 -246 2897 -212
rect 2841 -280 2897 -246
rect 2841 -314 2852 -280
rect 2886 -314 2897 -280
rect 2841 -348 2897 -314
rect 2841 -382 2852 -348
rect 2886 -382 2897 -348
rect 2841 -416 2897 -382
rect 2841 -450 2852 -416
rect 2886 -450 2897 -416
rect 2841 -484 2897 -450
rect 2841 -518 2852 -484
rect 2886 -518 2897 -484
rect 2841 -552 2897 -518
rect 2841 -586 2852 -552
rect 2886 -586 2897 -552
rect 2841 -620 2897 -586
rect 2841 -654 2852 -620
rect 2886 -654 2897 -620
rect 2841 -688 2897 -654
rect 2841 -722 2852 -688
rect 2886 -722 2897 -688
rect 2841 -756 2897 -722
rect 2841 -790 2852 -756
rect 2886 -790 2897 -756
rect 2841 -802 2897 -790
rect 3057 128 3113 198
rect 3057 94 3068 128
rect 3102 94 3113 128
rect 3057 60 3113 94
rect 3057 26 3068 60
rect 3102 26 3113 60
rect 3057 -8 3113 26
rect 3057 -42 3068 -8
rect 3102 -42 3113 -8
rect 3057 -76 3113 -42
rect 3057 -110 3068 -76
rect 3102 -110 3113 -76
rect 3057 -144 3113 -110
rect 3057 -178 3068 -144
rect 3102 -178 3113 -144
rect 3057 -212 3113 -178
rect 3057 -246 3068 -212
rect 3102 -246 3113 -212
rect 3057 -280 3113 -246
rect 3057 -314 3068 -280
rect 3102 -314 3113 -280
rect 3057 -348 3113 -314
rect 3057 -382 3068 -348
rect 3102 -382 3113 -348
rect 3057 -416 3113 -382
rect 3057 -450 3068 -416
rect 3102 -450 3113 -416
rect 3057 -484 3113 -450
rect 3057 -518 3068 -484
rect 3102 -518 3113 -484
rect 3057 -552 3113 -518
rect 3057 -586 3068 -552
rect 3102 -586 3113 -552
rect 3057 -620 3113 -586
rect 3057 -654 3068 -620
rect 3102 -654 3113 -620
rect 3057 -688 3113 -654
rect 3057 -722 3068 -688
rect 3102 -722 3113 -688
rect 3057 -756 3113 -722
rect 3057 -790 3068 -756
rect 3102 -790 3113 -756
rect 3057 -802 3113 -790
rect 3273 128 3326 198
rect 3273 94 3284 128
rect 3318 94 3326 128
rect 3273 60 3326 94
rect 3273 26 3284 60
rect 3318 26 3326 60
rect 3273 -8 3326 26
rect 3273 -42 3284 -8
rect 3318 -42 3326 -8
rect 3273 -76 3326 -42
rect 3273 -110 3284 -76
rect 3318 -110 3326 -76
rect 3273 -144 3326 -110
rect 3273 -178 3284 -144
rect 3318 -178 3326 -144
rect 3273 -212 3326 -178
rect 3273 -246 3284 -212
rect 3318 -246 3326 -212
rect 3273 -280 3326 -246
rect 3273 -314 3284 -280
rect 3318 -314 3326 -280
rect 3273 -348 3326 -314
rect 3273 -382 3284 -348
rect 3318 -382 3326 -348
rect 3273 -416 3326 -382
rect 3273 -450 3284 -416
rect 3318 -450 3326 -416
rect 3273 -484 3326 -450
rect 3273 -518 3284 -484
rect 3318 -518 3326 -484
rect 3273 -552 3326 -518
rect 3273 -586 3284 -552
rect 3318 -586 3326 -552
rect 3273 -620 3326 -586
rect 3273 -654 3284 -620
rect 3318 -654 3326 -620
rect 3273 -688 3326 -654
rect 3273 -722 3284 -688
rect 3318 -722 3326 -688
rect 3273 -756 3326 -722
rect 3273 -790 3284 -756
rect 3318 -790 3326 -756
rect 3273 -802 3326 -790
rect 3386 128 3439 198
rect 3386 94 3394 128
rect 3428 94 3439 128
rect 3386 60 3439 94
rect 3386 26 3394 60
rect 3428 26 3439 60
rect 3386 -8 3439 26
rect 3386 -42 3394 -8
rect 3428 -42 3439 -8
rect 3386 -76 3439 -42
rect 3386 -110 3394 -76
rect 3428 -110 3439 -76
rect 3386 -144 3439 -110
rect 3386 -178 3394 -144
rect 3428 -178 3439 -144
rect 3386 -212 3439 -178
rect 3386 -246 3394 -212
rect 3428 -246 3439 -212
rect 3386 -280 3439 -246
rect 3386 -314 3394 -280
rect 3428 -314 3439 -280
rect 3386 -348 3439 -314
rect 3386 -382 3394 -348
rect 3428 -382 3439 -348
rect 3386 -416 3439 -382
rect 3386 -450 3394 -416
rect 3428 -450 3439 -416
rect 3386 -484 3439 -450
rect 3386 -518 3394 -484
rect 3428 -518 3439 -484
rect 3386 -552 3439 -518
rect 3386 -586 3394 -552
rect 3428 -586 3439 -552
rect 3386 -620 3439 -586
rect 3386 -654 3394 -620
rect 3428 -654 3439 -620
rect 3386 -688 3439 -654
rect 3386 -722 3394 -688
rect 3428 -722 3439 -688
rect 3386 -756 3439 -722
rect 3386 -790 3394 -756
rect 3428 -790 3439 -756
rect 3386 -802 3439 -790
rect 3599 128 3652 198
rect 3599 94 3610 128
rect 3644 94 3652 128
rect 3599 60 3652 94
rect 3599 26 3610 60
rect 3644 26 3652 60
rect 3599 -8 3652 26
rect 3599 -42 3610 -8
rect 3644 -42 3652 -8
rect 3599 -76 3652 -42
rect 3599 -110 3610 -76
rect 3644 -110 3652 -76
rect 3599 -144 3652 -110
rect 3599 -178 3610 -144
rect 3644 -178 3652 -144
rect 3599 -212 3652 -178
rect 3599 -246 3610 -212
rect 3644 -246 3652 -212
rect 3599 -280 3652 -246
rect 3599 -314 3610 -280
rect 3644 -314 3652 -280
rect 3599 -348 3652 -314
rect 3599 -382 3610 -348
rect 3644 -382 3652 -348
rect 3599 -416 3652 -382
rect 3599 -450 3610 -416
rect 3644 -450 3652 -416
rect 3599 -484 3652 -450
rect 3599 -518 3610 -484
rect 3644 -518 3652 -484
rect 3599 -552 3652 -518
rect 3599 -586 3610 -552
rect 3644 -586 3652 -552
rect 3599 -620 3652 -586
rect 3599 -654 3610 -620
rect 3644 -654 3652 -620
rect 3599 -688 3652 -654
rect 3599 -722 3610 -688
rect 3644 -722 3652 -688
rect 3599 -756 3652 -722
rect 3599 -790 3610 -756
rect 3644 -790 3652 -756
rect 3599 -802 3652 -790
rect 3712 128 3765 198
rect 3712 94 3720 128
rect 3754 94 3765 128
rect 3712 60 3765 94
rect 3712 26 3720 60
rect 3754 26 3765 60
rect 3712 -8 3765 26
rect 3712 -42 3720 -8
rect 3754 -42 3765 -8
rect 3712 -76 3765 -42
rect 3712 -110 3720 -76
rect 3754 -110 3765 -76
rect 3712 -144 3765 -110
rect 3712 -178 3720 -144
rect 3754 -178 3765 -144
rect 3712 -212 3765 -178
rect 3712 -246 3720 -212
rect 3754 -246 3765 -212
rect 3712 -280 3765 -246
rect 3712 -314 3720 -280
rect 3754 -314 3765 -280
rect 3712 -348 3765 -314
rect 3712 -382 3720 -348
rect 3754 -382 3765 -348
rect 3712 -416 3765 -382
rect 3712 -450 3720 -416
rect 3754 -450 3765 -416
rect 3712 -484 3765 -450
rect 3712 -518 3720 -484
rect 3754 -518 3765 -484
rect 3712 -552 3765 -518
rect 3712 -586 3720 -552
rect 3754 -586 3765 -552
rect 3712 -620 3765 -586
rect 3712 -654 3720 -620
rect 3754 -654 3765 -620
rect 3712 -688 3765 -654
rect 3712 -722 3720 -688
rect 3754 -722 3765 -688
rect 3712 -756 3765 -722
rect 3712 -790 3720 -756
rect 3754 -790 3765 -756
rect 3712 -802 3765 -790
rect 3925 128 3978 198
rect 3925 94 3936 128
rect 3970 94 3978 128
rect 3925 60 3978 94
rect 3925 26 3936 60
rect 3970 26 3978 60
rect 3925 -8 3978 26
rect 3925 -42 3936 -8
rect 3970 -42 3978 -8
rect 3925 -76 3978 -42
rect 3925 -110 3936 -76
rect 3970 -110 3978 -76
rect 3925 -144 3978 -110
rect 3925 -178 3936 -144
rect 3970 -178 3978 -144
rect 3925 -212 3978 -178
rect 3925 -246 3936 -212
rect 3970 -246 3978 -212
rect 3925 -280 3978 -246
rect 3925 -314 3936 -280
rect 3970 -314 3978 -280
rect 3925 -348 3978 -314
rect 3925 -382 3936 -348
rect 3970 -382 3978 -348
rect 3925 -416 3978 -382
rect 3925 -450 3936 -416
rect 3970 -450 3978 -416
rect 3925 -484 3978 -450
rect 3925 -518 3936 -484
rect 3970 -518 3978 -484
rect 3925 -552 3978 -518
rect 3925 -586 3936 -552
rect 3970 -586 3978 -552
rect 3925 -620 3978 -586
rect 3925 -654 3936 -620
rect 3970 -654 3978 -620
rect 3925 -688 3978 -654
rect 3925 -722 3936 -688
rect 3970 -722 3978 -688
rect 3925 -756 3978 -722
rect 3925 -790 3936 -756
rect 3970 -790 3978 -756
rect 3925 -802 3978 -790
rect 4038 128 4091 198
rect 4038 94 4046 128
rect 4080 94 4091 128
rect 4038 60 4091 94
rect 4038 26 4046 60
rect 4080 26 4091 60
rect 4038 -8 4091 26
rect 4038 -42 4046 -8
rect 4080 -42 4091 -8
rect 4038 -76 4091 -42
rect 4038 -110 4046 -76
rect 4080 -110 4091 -76
rect 4038 -144 4091 -110
rect 4038 -178 4046 -144
rect 4080 -178 4091 -144
rect 4038 -212 4091 -178
rect 4038 -246 4046 -212
rect 4080 -246 4091 -212
rect 4038 -280 4091 -246
rect 4038 -314 4046 -280
rect 4080 -314 4091 -280
rect 4038 -348 4091 -314
rect 4038 -382 4046 -348
rect 4080 -382 4091 -348
rect 4038 -416 4091 -382
rect 4038 -450 4046 -416
rect 4080 -450 4091 -416
rect 4038 -484 4091 -450
rect 4038 -518 4046 -484
rect 4080 -518 4091 -484
rect 4038 -552 4091 -518
rect 4038 -586 4046 -552
rect 4080 -586 4091 -552
rect 4038 -620 4091 -586
rect 4038 -654 4046 -620
rect 4080 -654 4091 -620
rect 4038 -688 4091 -654
rect 4038 -722 4046 -688
rect 4080 -722 4091 -688
rect 4038 -756 4091 -722
rect 4038 -790 4046 -756
rect 4080 -790 4091 -756
rect 4038 -802 4091 -790
rect 4251 128 4304 198
rect 4251 94 4262 128
rect 4296 94 4304 128
rect 4251 60 4304 94
rect 4251 26 4262 60
rect 4296 26 4304 60
rect 4251 -8 4304 26
rect 4364 167 4372 201
rect 4406 167 4417 201
rect 4364 133 4417 167
rect 4364 99 4372 133
rect 4406 99 4417 133
rect 4364 65 4417 99
rect 4364 31 4372 65
rect 4406 31 4417 65
rect 4364 13 4417 31
rect 4577 201 4633 213
rect 4577 167 4588 201
rect 4622 167 4633 201
rect 4577 133 4633 167
rect 4577 99 4588 133
rect 4622 99 4633 133
rect 4577 65 4633 99
rect 4577 31 4588 65
rect 4622 31 4633 65
rect 4577 13 4633 31
rect 4793 201 4849 213
rect 4793 167 4804 201
rect 4838 167 4849 201
rect 4793 133 4849 167
rect 4793 99 4804 133
rect 4838 99 4849 133
rect 4793 65 4849 99
rect 4793 31 4804 65
rect 4838 31 4849 65
rect 4793 13 4849 31
rect 5009 201 5065 213
rect 5009 167 5020 201
rect 5054 167 5065 201
rect 5009 133 5065 167
rect 5009 99 5020 133
rect 5054 99 5065 133
rect 5009 65 5065 99
rect 5009 31 5020 65
rect 5054 31 5065 65
rect 5009 13 5065 31
rect 5225 201 5278 213
rect 5225 167 5236 201
rect 5270 167 5278 201
rect 5225 133 5278 167
rect 5225 99 5236 133
rect 5270 99 5278 133
rect 5225 65 5278 99
rect 5225 31 5236 65
rect 5270 31 5278 65
rect 5225 13 5278 31
rect 5354 128 5407 198
rect 5354 94 5362 128
rect 5396 94 5407 128
rect 5354 60 5407 94
rect 5354 26 5362 60
rect 5396 26 5407 60
rect 4251 -42 4262 -8
rect 4296 -42 4304 -8
rect 5354 -8 5407 26
rect 4251 -76 4304 -42
rect 4251 -110 4262 -76
rect 4296 -110 4304 -76
rect 5354 -42 5362 -8
rect 5396 -42 5407 -8
rect 5354 -76 5407 -42
rect 4251 -144 4304 -110
rect 4251 -178 4262 -144
rect 4296 -178 4304 -144
rect 4251 -212 4304 -178
rect 5354 -110 5362 -76
rect 5396 -110 5407 -76
rect 5354 -144 5407 -110
rect 5354 -178 5362 -144
rect 5396 -178 5407 -144
rect 4251 -246 4262 -212
rect 4296 -246 4304 -212
rect 4251 -280 4304 -246
rect 4251 -314 4262 -280
rect 4296 -314 4304 -280
rect 4251 -348 4304 -314
rect 4251 -382 4262 -348
rect 4296 -382 4304 -348
rect 4251 -416 4304 -382
rect 4251 -450 4262 -416
rect 4296 -450 4304 -416
rect 4251 -484 4304 -450
rect 4251 -518 4262 -484
rect 4296 -518 4304 -484
rect 4251 -552 4304 -518
rect 4251 -586 4262 -552
rect 4296 -586 4304 -552
rect 4251 -620 4304 -586
rect 4251 -654 4262 -620
rect 4296 -654 4304 -620
rect 4251 -688 4304 -654
rect 4251 -722 4262 -688
rect 4296 -722 4304 -688
rect 4251 -756 4304 -722
rect 4251 -790 4262 -756
rect 4296 -790 4304 -756
rect 4251 -802 4304 -790
rect 4364 -280 4417 -202
rect 4364 -314 4372 -280
rect 4406 -314 4417 -280
rect 4364 -348 4417 -314
rect 4364 -382 4372 -348
rect 4406 -382 4417 -348
rect 4364 -416 4417 -382
rect 4364 -450 4372 -416
rect 4406 -450 4417 -416
rect 4364 -484 4417 -450
rect 4364 -518 4372 -484
rect 4406 -518 4417 -484
rect 4364 -552 4417 -518
rect 4364 -586 4372 -552
rect 4406 -586 4417 -552
rect 4364 -620 4417 -586
rect 4364 -654 4372 -620
rect 4406 -654 4417 -620
rect 4364 -688 4417 -654
rect 4364 -722 4372 -688
rect 4406 -722 4417 -688
rect 4364 -756 4417 -722
rect 4364 -790 4372 -756
rect 4406 -790 4417 -756
rect 4364 -802 4417 -790
rect 4617 -280 4673 -202
rect 4617 -314 4628 -280
rect 4662 -314 4673 -280
rect 4617 -348 4673 -314
rect 4617 -382 4628 -348
rect 4662 -382 4673 -348
rect 4617 -416 4673 -382
rect 4617 -450 4628 -416
rect 4662 -450 4673 -416
rect 4617 -484 4673 -450
rect 4617 -518 4628 -484
rect 4662 -518 4673 -484
rect 4617 -552 4673 -518
rect 4617 -586 4628 -552
rect 4662 -586 4673 -552
rect 4617 -620 4673 -586
rect 4617 -654 4628 -620
rect 4662 -654 4673 -620
rect 4617 -688 4673 -654
rect 4617 -722 4628 -688
rect 4662 -722 4673 -688
rect 4617 -756 4673 -722
rect 4617 -790 4628 -756
rect 4662 -790 4673 -756
rect 4617 -802 4673 -790
rect 4773 -280 4829 -202
rect 4773 -314 4784 -280
rect 4818 -314 4829 -280
rect 4773 -348 4829 -314
rect 4773 -382 4784 -348
rect 4818 -382 4829 -348
rect 4773 -416 4829 -382
rect 4773 -450 4784 -416
rect 4818 -450 4829 -416
rect 4773 -484 4829 -450
rect 4773 -518 4784 -484
rect 4818 -518 4829 -484
rect 4773 -552 4829 -518
rect 4773 -586 4784 -552
rect 4818 -586 4829 -552
rect 4773 -620 4829 -586
rect 4773 -654 4784 -620
rect 4818 -654 4829 -620
rect 4773 -688 4829 -654
rect 4773 -722 4784 -688
rect 4818 -722 4829 -688
rect 4773 -756 4829 -722
rect 4773 -790 4784 -756
rect 4818 -790 4829 -756
rect 4773 -802 4829 -790
rect 4929 -280 4985 -202
rect 4929 -314 4940 -280
rect 4974 -314 4985 -280
rect 4929 -348 4985 -314
rect 4929 -382 4940 -348
rect 4974 -382 4985 -348
rect 4929 -416 4985 -382
rect 4929 -450 4940 -416
rect 4974 -450 4985 -416
rect 4929 -484 4985 -450
rect 4929 -518 4940 -484
rect 4974 -518 4985 -484
rect 4929 -552 4985 -518
rect 4929 -586 4940 -552
rect 4974 -586 4985 -552
rect 4929 -620 4985 -586
rect 4929 -654 4940 -620
rect 4974 -654 4985 -620
rect 4929 -688 4985 -654
rect 4929 -722 4940 -688
rect 4974 -722 4985 -688
rect 4929 -756 4985 -722
rect 4929 -790 4940 -756
rect 4974 -790 4985 -756
rect 4929 -802 4985 -790
rect 5085 -280 5141 -202
rect 5085 -314 5096 -280
rect 5130 -314 5141 -280
rect 5085 -348 5141 -314
rect 5085 -382 5096 -348
rect 5130 -382 5141 -348
rect 5085 -416 5141 -382
rect 5085 -450 5096 -416
rect 5130 -450 5141 -416
rect 5085 -484 5141 -450
rect 5085 -518 5096 -484
rect 5130 -518 5141 -484
rect 5085 -552 5141 -518
rect 5085 -586 5096 -552
rect 5130 -586 5141 -552
rect 5085 -620 5141 -586
rect 5085 -654 5096 -620
rect 5130 -654 5141 -620
rect 5085 -688 5141 -654
rect 5085 -722 5096 -688
rect 5130 -722 5141 -688
rect 5085 -756 5141 -722
rect 5085 -790 5096 -756
rect 5130 -790 5141 -756
rect 5085 -802 5141 -790
rect 5241 -280 5294 -202
rect 5241 -314 5252 -280
rect 5286 -314 5294 -280
rect 5241 -348 5294 -314
rect 5241 -382 5252 -348
rect 5286 -382 5294 -348
rect 5241 -416 5294 -382
rect 5241 -450 5252 -416
rect 5286 -450 5294 -416
rect 5241 -484 5294 -450
rect 5241 -518 5252 -484
rect 5286 -518 5294 -484
rect 5241 -552 5294 -518
rect 5241 -586 5252 -552
rect 5286 -586 5294 -552
rect 5241 -620 5294 -586
rect 5241 -654 5252 -620
rect 5286 -654 5294 -620
rect 5241 -688 5294 -654
rect 5241 -722 5252 -688
rect 5286 -722 5294 -688
rect 5241 -756 5294 -722
rect 5241 -790 5252 -756
rect 5286 -790 5294 -756
rect 5241 -802 5294 -790
rect 5354 -212 5407 -178
rect 5354 -246 5362 -212
rect 5396 -246 5407 -212
rect 5354 -280 5407 -246
rect 5354 -314 5362 -280
rect 5396 -314 5407 -280
rect 5354 -348 5407 -314
rect 5354 -382 5362 -348
rect 5396 -382 5407 -348
rect 5354 -416 5407 -382
rect 5354 -450 5362 -416
rect 5396 -450 5407 -416
rect 5354 -484 5407 -450
rect 5354 -518 5362 -484
rect 5396 -518 5407 -484
rect 5354 -552 5407 -518
rect 5354 -586 5362 -552
rect 5396 -586 5407 -552
rect 5354 -620 5407 -586
rect 5354 -654 5362 -620
rect 5396 -654 5407 -620
rect 5354 -688 5407 -654
rect 5354 -722 5362 -688
rect 5396 -722 5407 -688
rect 5354 -756 5407 -722
rect 5354 -790 5362 -756
rect 5396 -790 5407 -756
rect 5354 -802 5407 -790
rect 5507 128 5563 198
rect 5507 94 5518 128
rect 5552 94 5563 128
rect 5507 60 5563 94
rect 5507 26 5518 60
rect 5552 26 5563 60
rect 5507 -8 5563 26
rect 5507 -42 5518 -8
rect 5552 -42 5563 -8
rect 5507 -76 5563 -42
rect 5507 -110 5518 -76
rect 5552 -110 5563 -76
rect 5507 -144 5563 -110
rect 5507 -178 5518 -144
rect 5552 -178 5563 -144
rect 5507 -212 5563 -178
rect 5507 -246 5518 -212
rect 5552 -246 5563 -212
rect 5507 -280 5563 -246
rect 5507 -314 5518 -280
rect 5552 -314 5563 -280
rect 5507 -348 5563 -314
rect 5507 -382 5518 -348
rect 5552 -382 5563 -348
rect 5507 -416 5563 -382
rect 5507 -450 5518 -416
rect 5552 -450 5563 -416
rect 5507 -484 5563 -450
rect 5507 -518 5518 -484
rect 5552 -518 5563 -484
rect 5507 -552 5563 -518
rect 5507 -586 5518 -552
rect 5552 -586 5563 -552
rect 5507 -620 5563 -586
rect 5507 -654 5518 -620
rect 5552 -654 5563 -620
rect 5507 -688 5563 -654
rect 5507 -722 5518 -688
rect 5552 -722 5563 -688
rect 5507 -756 5563 -722
rect 5507 -790 5518 -756
rect 5552 -790 5563 -756
rect 5507 -802 5563 -790
rect 5663 128 5716 198
rect 5663 94 5674 128
rect 5708 94 5716 128
rect 5663 60 5716 94
rect 5663 26 5674 60
rect 5708 26 5716 60
rect 5663 -8 5716 26
rect 5663 -42 5674 -8
rect 5708 -42 5716 -8
rect 5663 -76 5716 -42
rect 5663 -110 5674 -76
rect 5708 -110 5716 -76
rect 5663 -144 5716 -110
rect 5663 -178 5674 -144
rect 5708 -178 5716 -144
rect 5663 -212 5716 -178
rect 5663 -246 5674 -212
rect 5708 -246 5716 -212
rect 5663 -280 5716 -246
rect 5663 -314 5674 -280
rect 5708 -314 5716 -280
rect 5663 -348 5716 -314
rect 5663 -382 5674 -348
rect 5708 -382 5716 -348
rect 5663 -416 5716 -382
rect 5663 -450 5674 -416
rect 5708 -450 5716 -416
rect 5663 -484 5716 -450
rect 5663 -518 5674 -484
rect 5708 -518 5716 -484
rect 5663 -552 5716 -518
rect 5663 -586 5674 -552
rect 5708 -586 5716 -552
rect 5663 -620 5716 -586
rect 5663 -654 5674 -620
rect 5708 -654 5716 -620
rect 5663 -688 5716 -654
rect 5663 -722 5674 -688
rect 5708 -722 5716 -688
rect 5663 -756 5716 -722
rect 5663 -790 5674 -756
rect 5708 -790 5716 -756
rect 5663 -802 5716 -790
<< mvpdiff >>
rect 66 2795 119 2865
rect 66 2761 74 2795
rect 108 2761 119 2795
rect 66 2727 119 2761
rect 66 2693 74 2727
rect 108 2693 119 2727
rect 66 2659 119 2693
rect 66 2625 74 2659
rect 108 2625 119 2659
rect 66 2591 119 2625
rect 66 2557 74 2591
rect 108 2557 119 2591
rect 66 2523 119 2557
rect 66 2489 74 2523
rect 108 2489 119 2523
rect 66 2455 119 2489
rect 66 2421 74 2455
rect 108 2421 119 2455
rect 66 2387 119 2421
rect 66 2353 74 2387
rect 108 2353 119 2387
rect 66 2319 119 2353
rect 66 2285 74 2319
rect 108 2285 119 2319
rect 66 2251 119 2285
rect 66 2217 74 2251
rect 108 2217 119 2251
rect 66 2183 119 2217
rect 66 2149 74 2183
rect 108 2149 119 2183
rect 66 2115 119 2149
rect 66 2081 74 2115
rect 108 2081 119 2115
rect 66 2047 119 2081
rect 66 2013 74 2047
rect 108 2013 119 2047
rect 66 1979 119 2013
rect 66 1945 74 1979
rect 108 1945 119 1979
rect 66 1911 119 1945
rect 66 1877 74 1911
rect 108 1877 119 1911
rect 66 1865 119 1877
rect 219 2795 275 2865
rect 219 2761 230 2795
rect 264 2761 275 2795
rect 219 2727 275 2761
rect 219 2693 230 2727
rect 264 2693 275 2727
rect 219 2659 275 2693
rect 219 2625 230 2659
rect 264 2625 275 2659
rect 219 2591 275 2625
rect 219 2557 230 2591
rect 264 2557 275 2591
rect 219 2523 275 2557
rect 219 2489 230 2523
rect 264 2489 275 2523
rect 219 2455 275 2489
rect 219 2421 230 2455
rect 264 2421 275 2455
rect 219 2387 275 2421
rect 219 2353 230 2387
rect 264 2353 275 2387
rect 219 2319 275 2353
rect 219 2285 230 2319
rect 264 2285 275 2319
rect 219 2251 275 2285
rect 219 2217 230 2251
rect 264 2217 275 2251
rect 219 2183 275 2217
rect 219 2149 230 2183
rect 264 2149 275 2183
rect 219 2115 275 2149
rect 219 2081 230 2115
rect 264 2081 275 2115
rect 219 2047 275 2081
rect 219 2013 230 2047
rect 264 2013 275 2047
rect 219 1979 275 2013
rect 219 1945 230 1979
rect 264 1945 275 1979
rect 219 1911 275 1945
rect 219 1877 230 1911
rect 264 1877 275 1911
rect 219 1865 275 1877
rect 375 2795 428 2865
rect 375 2761 386 2795
rect 420 2761 428 2795
rect 375 2727 428 2761
rect 375 2693 386 2727
rect 420 2693 428 2727
rect 375 2659 428 2693
rect 375 2625 386 2659
rect 420 2625 428 2659
rect 375 2591 428 2625
rect 375 2557 386 2591
rect 420 2557 428 2591
rect 375 2523 428 2557
rect 375 2489 386 2523
rect 420 2489 428 2523
rect 375 2455 428 2489
rect 375 2421 386 2455
rect 420 2421 428 2455
rect 375 2387 428 2421
rect 375 2353 386 2387
rect 420 2353 428 2387
rect 375 2319 428 2353
rect 375 2285 386 2319
rect 420 2285 428 2319
rect 375 2251 428 2285
rect 375 2217 386 2251
rect 420 2217 428 2251
rect 375 2183 428 2217
rect 375 2149 386 2183
rect 420 2149 428 2183
rect 375 2115 428 2149
rect 375 2081 386 2115
rect 420 2081 428 2115
rect 375 2047 428 2081
rect 375 2013 386 2047
rect 420 2013 428 2047
rect 375 1979 428 2013
rect 375 1945 386 1979
rect 420 1945 428 1979
rect 375 1911 428 1945
rect 375 1877 386 1911
rect 420 1877 428 1911
rect 375 1865 428 1877
rect 488 2795 541 2865
rect 488 2761 496 2795
rect 530 2761 541 2795
rect 488 2727 541 2761
rect 488 2693 496 2727
rect 530 2693 541 2727
rect 488 2659 541 2693
rect 488 2625 496 2659
rect 530 2625 541 2659
rect 488 2591 541 2625
rect 488 2557 496 2591
rect 530 2557 541 2591
rect 488 2523 541 2557
rect 488 2489 496 2523
rect 530 2489 541 2523
rect 488 2455 541 2489
rect 488 2421 496 2455
rect 530 2421 541 2455
rect 488 2387 541 2421
rect 488 2353 496 2387
rect 530 2353 541 2387
rect 488 2319 541 2353
rect 488 2285 496 2319
rect 530 2285 541 2319
rect 488 2251 541 2285
rect 488 2217 496 2251
rect 530 2217 541 2251
rect 488 2183 541 2217
rect 488 2149 496 2183
rect 530 2149 541 2183
rect 488 2115 541 2149
rect 488 2081 496 2115
rect 530 2081 541 2115
rect 488 2047 541 2081
rect 488 2013 496 2047
rect 530 2013 541 2047
rect 488 1979 541 2013
rect 488 1945 496 1979
rect 530 1945 541 1979
rect 488 1911 541 1945
rect 488 1877 496 1911
rect 530 1877 541 1911
rect 488 1865 541 1877
rect 701 2795 757 2865
rect 701 2761 712 2795
rect 746 2761 757 2795
rect 701 2727 757 2761
rect 701 2693 712 2727
rect 746 2693 757 2727
rect 701 2659 757 2693
rect 701 2625 712 2659
rect 746 2625 757 2659
rect 701 2591 757 2625
rect 701 2557 712 2591
rect 746 2557 757 2591
rect 701 2523 757 2557
rect 701 2489 712 2523
rect 746 2489 757 2523
rect 701 2455 757 2489
rect 701 2421 712 2455
rect 746 2421 757 2455
rect 701 2387 757 2421
rect 701 2353 712 2387
rect 746 2353 757 2387
rect 701 2319 757 2353
rect 701 2285 712 2319
rect 746 2285 757 2319
rect 701 2251 757 2285
rect 701 2217 712 2251
rect 746 2217 757 2251
rect 701 2183 757 2217
rect 701 2149 712 2183
rect 746 2149 757 2183
rect 701 2115 757 2149
rect 701 2081 712 2115
rect 746 2081 757 2115
rect 701 2047 757 2081
rect 701 2013 712 2047
rect 746 2013 757 2047
rect 701 1979 757 2013
rect 701 1945 712 1979
rect 746 1945 757 1979
rect 701 1911 757 1945
rect 701 1877 712 1911
rect 746 1877 757 1911
rect 701 1865 757 1877
rect 917 2795 973 2865
rect 917 2761 928 2795
rect 962 2761 973 2795
rect 917 2727 973 2761
rect 917 2693 928 2727
rect 962 2693 973 2727
rect 917 2659 973 2693
rect 917 2625 928 2659
rect 962 2625 973 2659
rect 917 2591 973 2625
rect 917 2557 928 2591
rect 962 2557 973 2591
rect 917 2523 973 2557
rect 917 2489 928 2523
rect 962 2489 973 2523
rect 917 2455 973 2489
rect 917 2421 928 2455
rect 962 2421 973 2455
rect 917 2387 973 2421
rect 917 2353 928 2387
rect 962 2353 973 2387
rect 917 2319 973 2353
rect 917 2285 928 2319
rect 962 2285 973 2319
rect 917 2251 973 2285
rect 917 2217 928 2251
rect 962 2217 973 2251
rect 917 2183 973 2217
rect 917 2149 928 2183
rect 962 2149 973 2183
rect 917 2115 973 2149
rect 917 2081 928 2115
rect 962 2081 973 2115
rect 917 2047 973 2081
rect 917 2013 928 2047
rect 962 2013 973 2047
rect 917 1979 973 2013
rect 917 1945 928 1979
rect 962 1945 973 1979
rect 917 1911 973 1945
rect 917 1877 928 1911
rect 962 1877 973 1911
rect 917 1865 973 1877
rect 1073 2795 1129 2865
rect 1073 2761 1084 2795
rect 1118 2761 1129 2795
rect 1073 2727 1129 2761
rect 1073 2693 1084 2727
rect 1118 2693 1129 2727
rect 1073 2659 1129 2693
rect 1073 2625 1084 2659
rect 1118 2625 1129 2659
rect 1073 2591 1129 2625
rect 1073 2557 1084 2591
rect 1118 2557 1129 2591
rect 1073 2523 1129 2557
rect 1073 2489 1084 2523
rect 1118 2489 1129 2523
rect 1073 2455 1129 2489
rect 1073 2421 1084 2455
rect 1118 2421 1129 2455
rect 1073 2387 1129 2421
rect 1073 2353 1084 2387
rect 1118 2353 1129 2387
rect 1073 2319 1129 2353
rect 1073 2285 1084 2319
rect 1118 2285 1129 2319
rect 1073 2251 1129 2285
rect 1073 2217 1084 2251
rect 1118 2217 1129 2251
rect 1073 2183 1129 2217
rect 1073 2149 1084 2183
rect 1118 2149 1129 2183
rect 1073 2115 1129 2149
rect 1073 2081 1084 2115
rect 1118 2081 1129 2115
rect 1073 2047 1129 2081
rect 1073 2013 1084 2047
rect 1118 2013 1129 2047
rect 1073 1979 1129 2013
rect 1073 1945 1084 1979
rect 1118 1945 1129 1979
rect 1073 1911 1129 1945
rect 1073 1877 1084 1911
rect 1118 1877 1129 1911
rect 1073 1865 1129 1877
rect 1229 2795 1282 2865
rect 1229 2761 1240 2795
rect 1274 2761 1282 2795
rect 1229 2727 1282 2761
rect 1229 2693 1240 2727
rect 1274 2693 1282 2727
rect 1229 2659 1282 2693
rect 1229 2625 1240 2659
rect 1274 2625 1282 2659
rect 1229 2591 1282 2625
rect 1229 2557 1240 2591
rect 1274 2557 1282 2591
rect 1229 2523 1282 2557
rect 1229 2489 1240 2523
rect 1274 2489 1282 2523
rect 1229 2455 1282 2489
rect 1229 2421 1240 2455
rect 1274 2421 1282 2455
rect 1229 2387 1282 2421
rect 1229 2353 1240 2387
rect 1274 2353 1282 2387
rect 1229 2319 1282 2353
rect 1229 2285 1240 2319
rect 1274 2285 1282 2319
rect 1229 2251 1282 2285
rect 1229 2217 1240 2251
rect 1274 2217 1282 2251
rect 1229 2183 1282 2217
rect 1229 2149 1240 2183
rect 1274 2149 1282 2183
rect 1229 2115 1282 2149
rect 1229 2081 1240 2115
rect 1274 2081 1282 2115
rect 1229 2047 1282 2081
rect 1229 2013 1240 2047
rect 1274 2013 1282 2047
rect 1229 1979 1282 2013
rect 1229 1945 1240 1979
rect 1274 1945 1282 1979
rect 1229 1911 1282 1945
rect 1229 1877 1240 1911
rect 1274 1877 1282 1911
rect 1229 1865 1282 1877
rect 1392 2795 1445 2865
rect 1392 2761 1400 2795
rect 1434 2761 1445 2795
rect 1392 2727 1445 2761
rect 1392 2693 1400 2727
rect 1434 2693 1445 2727
rect 1392 2659 1445 2693
rect 1392 2625 1400 2659
rect 1434 2625 1445 2659
rect 1392 2591 1445 2625
rect 1392 2557 1400 2591
rect 1434 2557 1445 2591
rect 1392 2523 1445 2557
rect 1392 2489 1400 2523
rect 1434 2489 1445 2523
rect 1392 2455 1445 2489
rect 1392 2421 1400 2455
rect 1434 2421 1445 2455
rect 1392 2387 1445 2421
rect 1392 2353 1400 2387
rect 1434 2353 1445 2387
rect 1392 2319 1445 2353
rect 1392 2285 1400 2319
rect 1434 2285 1445 2319
rect 1392 2251 1445 2285
rect 1392 2217 1400 2251
rect 1434 2217 1445 2251
rect 1392 2183 1445 2217
rect 1392 2149 1400 2183
rect 1434 2149 1445 2183
rect 1392 2115 1445 2149
rect 1392 2081 1400 2115
rect 1434 2081 1445 2115
rect 1392 2047 1445 2081
rect 1392 2013 1400 2047
rect 1434 2013 1445 2047
rect 1392 1979 1445 2013
rect 1392 1945 1400 1979
rect 1434 1945 1445 1979
rect 1392 1911 1445 1945
rect 1392 1877 1400 1911
rect 1434 1877 1445 1911
rect 1392 1865 1445 1877
rect 1605 2795 1661 2865
rect 1605 2761 1616 2795
rect 1650 2761 1661 2795
rect 1605 2727 1661 2761
rect 1605 2693 1616 2727
rect 1650 2693 1661 2727
rect 1605 2659 1661 2693
rect 1605 2625 1616 2659
rect 1650 2625 1661 2659
rect 1605 2591 1661 2625
rect 1605 2557 1616 2591
rect 1650 2557 1661 2591
rect 1605 2523 1661 2557
rect 1605 2489 1616 2523
rect 1650 2489 1661 2523
rect 1605 2455 1661 2489
rect 1605 2421 1616 2455
rect 1650 2421 1661 2455
rect 1605 2387 1661 2421
rect 1605 2353 1616 2387
rect 1650 2353 1661 2387
rect 1605 2319 1661 2353
rect 1605 2285 1616 2319
rect 1650 2285 1661 2319
rect 1605 2251 1661 2285
rect 1605 2217 1616 2251
rect 1650 2217 1661 2251
rect 1605 2183 1661 2217
rect 1605 2149 1616 2183
rect 1650 2149 1661 2183
rect 1605 2115 1661 2149
rect 1605 2081 1616 2115
rect 1650 2081 1661 2115
rect 1605 2047 1661 2081
rect 1605 2013 1616 2047
rect 1650 2013 1661 2047
rect 1605 1979 1661 2013
rect 1605 1945 1616 1979
rect 1650 1945 1661 1979
rect 1605 1911 1661 1945
rect 1605 1877 1616 1911
rect 1650 1877 1661 1911
rect 1605 1865 1661 1877
rect 1761 2795 1817 2865
rect 1761 2761 1772 2795
rect 1806 2761 1817 2795
rect 1761 2727 1817 2761
rect 1761 2693 1772 2727
rect 1806 2693 1817 2727
rect 1761 2659 1817 2693
rect 1761 2625 1772 2659
rect 1806 2625 1817 2659
rect 1761 2591 1817 2625
rect 1761 2557 1772 2591
rect 1806 2557 1817 2591
rect 1761 2523 1817 2557
rect 1761 2489 1772 2523
rect 1806 2489 1817 2523
rect 1761 2455 1817 2489
rect 1761 2421 1772 2455
rect 1806 2421 1817 2455
rect 1761 2387 1817 2421
rect 1761 2353 1772 2387
rect 1806 2353 1817 2387
rect 1761 2319 1817 2353
rect 1761 2285 1772 2319
rect 1806 2285 1817 2319
rect 1761 2251 1817 2285
rect 1761 2217 1772 2251
rect 1806 2217 1817 2251
rect 1761 2183 1817 2217
rect 1761 2149 1772 2183
rect 1806 2149 1817 2183
rect 1761 2115 1817 2149
rect 1761 2081 1772 2115
rect 1806 2081 1817 2115
rect 1761 2047 1817 2081
rect 1761 2013 1772 2047
rect 1806 2013 1817 2047
rect 1761 1979 1817 2013
rect 1761 1945 1772 1979
rect 1806 1945 1817 1979
rect 1761 1911 1817 1945
rect 1761 1877 1772 1911
rect 1806 1877 1817 1911
rect 1761 1865 1817 1877
rect 1917 2795 1973 2865
rect 1917 2761 1928 2795
rect 1962 2761 1973 2795
rect 1917 2727 1973 2761
rect 1917 2693 1928 2727
rect 1962 2693 1973 2727
rect 1917 2659 1973 2693
rect 1917 2625 1928 2659
rect 1962 2625 1973 2659
rect 1917 2591 1973 2625
rect 1917 2557 1928 2591
rect 1962 2557 1973 2591
rect 1917 2523 1973 2557
rect 1917 2489 1928 2523
rect 1962 2489 1973 2523
rect 1917 2455 1973 2489
rect 1917 2421 1928 2455
rect 1962 2421 1973 2455
rect 1917 2387 1973 2421
rect 1917 2353 1928 2387
rect 1962 2353 1973 2387
rect 1917 2319 1973 2353
rect 1917 2285 1928 2319
rect 1962 2285 1973 2319
rect 1917 2251 1973 2285
rect 1917 2217 1928 2251
rect 1962 2217 1973 2251
rect 1917 2183 1973 2217
rect 1917 2149 1928 2183
rect 1962 2149 1973 2183
rect 1917 2115 1973 2149
rect 1917 2081 1928 2115
rect 1962 2081 1973 2115
rect 1917 2047 1973 2081
rect 1917 2013 1928 2047
rect 1962 2013 1973 2047
rect 1917 1979 1973 2013
rect 1917 1945 1928 1979
rect 1962 1945 1973 1979
rect 1917 1911 1973 1945
rect 1917 1877 1928 1911
rect 1962 1877 1973 1911
rect 1917 1865 1973 1877
rect 2073 2795 2129 2865
rect 2073 2761 2084 2795
rect 2118 2761 2129 2795
rect 2073 2727 2129 2761
rect 2073 2693 2084 2727
rect 2118 2693 2129 2727
rect 2073 2659 2129 2693
rect 2073 2625 2084 2659
rect 2118 2625 2129 2659
rect 2073 2591 2129 2625
rect 2073 2557 2084 2591
rect 2118 2557 2129 2591
rect 2073 2523 2129 2557
rect 2073 2489 2084 2523
rect 2118 2489 2129 2523
rect 2073 2455 2129 2489
rect 2073 2421 2084 2455
rect 2118 2421 2129 2455
rect 2073 2387 2129 2421
rect 2073 2353 2084 2387
rect 2118 2353 2129 2387
rect 2073 2319 2129 2353
rect 2073 2285 2084 2319
rect 2118 2285 2129 2319
rect 2073 2251 2129 2285
rect 2073 2217 2084 2251
rect 2118 2217 2129 2251
rect 2073 2183 2129 2217
rect 2073 2149 2084 2183
rect 2118 2149 2129 2183
rect 2073 2115 2129 2149
rect 2073 2081 2084 2115
rect 2118 2081 2129 2115
rect 2073 2047 2129 2081
rect 2073 2013 2084 2047
rect 2118 2013 2129 2047
rect 2073 1979 2129 2013
rect 2073 1945 2084 1979
rect 2118 1945 2129 1979
rect 2073 1911 2129 1945
rect 2073 1877 2084 1911
rect 2118 1877 2129 1911
rect 2073 1865 2129 1877
rect 2229 2795 2285 2865
rect 2229 2761 2240 2795
rect 2274 2761 2285 2795
rect 2229 2727 2285 2761
rect 2229 2693 2240 2727
rect 2274 2693 2285 2727
rect 2229 2659 2285 2693
rect 2229 2625 2240 2659
rect 2274 2625 2285 2659
rect 2229 2591 2285 2625
rect 2229 2557 2240 2591
rect 2274 2557 2285 2591
rect 2229 2523 2285 2557
rect 2229 2489 2240 2523
rect 2274 2489 2285 2523
rect 2229 2455 2285 2489
rect 2229 2421 2240 2455
rect 2274 2421 2285 2455
rect 2229 2387 2285 2421
rect 2229 2353 2240 2387
rect 2274 2353 2285 2387
rect 2229 2319 2285 2353
rect 2229 2285 2240 2319
rect 2274 2285 2285 2319
rect 2229 2251 2285 2285
rect 2229 2217 2240 2251
rect 2274 2217 2285 2251
rect 2229 2183 2285 2217
rect 2229 2149 2240 2183
rect 2274 2149 2285 2183
rect 2229 2115 2285 2149
rect 2229 2081 2240 2115
rect 2274 2081 2285 2115
rect 2229 2047 2285 2081
rect 2229 2013 2240 2047
rect 2274 2013 2285 2047
rect 2229 1979 2285 2013
rect 2229 1945 2240 1979
rect 2274 1945 2285 1979
rect 2229 1911 2285 1945
rect 2229 1877 2240 1911
rect 2274 1877 2285 1911
rect 2229 1865 2285 1877
rect 2385 2795 2438 2865
rect 2385 2761 2396 2795
rect 2430 2761 2438 2795
rect 2385 2727 2438 2761
rect 2385 2693 2396 2727
rect 2430 2693 2438 2727
rect 2385 2659 2438 2693
rect 2385 2625 2396 2659
rect 2430 2625 2438 2659
rect 2385 2591 2438 2625
rect 2385 2557 2396 2591
rect 2430 2557 2438 2591
rect 2385 2523 2438 2557
rect 2385 2489 2396 2523
rect 2430 2489 2438 2523
rect 2764 2795 2817 2865
rect 2764 2761 2772 2795
rect 2806 2761 2817 2795
rect 2764 2727 2817 2761
rect 2764 2693 2772 2727
rect 2806 2693 2817 2727
rect 2764 2659 2817 2693
rect 2764 2625 2772 2659
rect 2806 2625 2817 2659
rect 2764 2591 2817 2625
rect 2764 2557 2772 2591
rect 2806 2557 2817 2591
rect 2764 2523 2817 2557
rect 2385 2455 2438 2489
rect 2764 2489 2772 2523
rect 2806 2489 2817 2523
rect 2385 2421 2396 2455
rect 2430 2421 2438 2455
rect 2385 2387 2438 2421
rect 2385 2353 2396 2387
rect 2430 2353 2438 2387
rect 2385 2319 2438 2353
rect 2385 2285 2396 2319
rect 2430 2285 2438 2319
rect 2385 2251 2438 2285
rect 2385 2217 2396 2251
rect 2430 2217 2438 2251
rect 2385 2183 2438 2217
rect 2385 2149 2396 2183
rect 2430 2149 2438 2183
rect 2385 2115 2438 2149
rect 2385 2081 2396 2115
rect 2430 2081 2438 2115
rect 2385 2047 2438 2081
rect 2385 2013 2396 2047
rect 2430 2013 2438 2047
rect 2385 1979 2438 2013
rect 2385 1945 2396 1979
rect 2430 1945 2438 1979
rect 2385 1911 2438 1945
rect 2385 1877 2396 1911
rect 2430 1877 2438 1911
rect 2385 1865 2438 1877
rect 2498 2387 2551 2465
rect 2498 2353 2506 2387
rect 2540 2353 2551 2387
rect 2498 2319 2551 2353
rect 2498 2285 2506 2319
rect 2540 2285 2551 2319
rect 2498 2251 2551 2285
rect 2498 2217 2506 2251
rect 2540 2217 2551 2251
rect 2498 2183 2551 2217
rect 2498 2149 2506 2183
rect 2540 2149 2551 2183
rect 2498 2115 2551 2149
rect 2498 2081 2506 2115
rect 2540 2081 2551 2115
rect 2498 2047 2551 2081
rect 2498 2013 2506 2047
rect 2540 2013 2551 2047
rect 2498 1979 2551 2013
rect 2498 1945 2506 1979
rect 2540 1945 2551 1979
rect 2498 1911 2551 1945
rect 2498 1877 2506 1911
rect 2540 1877 2551 1911
rect 2498 1865 2551 1877
rect 2651 2387 2704 2465
rect 2651 2353 2662 2387
rect 2696 2353 2704 2387
rect 2651 2319 2704 2353
rect 2651 2285 2662 2319
rect 2696 2285 2704 2319
rect 2651 2251 2704 2285
rect 2651 2217 2662 2251
rect 2696 2217 2704 2251
rect 2651 2183 2704 2217
rect 2651 2149 2662 2183
rect 2696 2149 2704 2183
rect 2651 2115 2704 2149
rect 2651 2081 2662 2115
rect 2696 2081 2704 2115
rect 2651 2047 2704 2081
rect 2651 2013 2662 2047
rect 2696 2013 2704 2047
rect 2651 1979 2704 2013
rect 2651 1945 2662 1979
rect 2696 1945 2704 1979
rect 2651 1911 2704 1945
rect 2651 1877 2662 1911
rect 2696 1877 2704 1911
rect 2651 1865 2704 1877
rect 2764 2455 2817 2489
rect 2764 2421 2772 2455
rect 2806 2421 2817 2455
rect 2764 2387 2817 2421
rect 2764 2353 2772 2387
rect 2806 2353 2817 2387
rect 2764 2319 2817 2353
rect 2764 2285 2772 2319
rect 2806 2285 2817 2319
rect 2764 2251 2817 2285
rect 2764 2217 2772 2251
rect 2806 2217 2817 2251
rect 2764 2183 2817 2217
rect 2764 2149 2772 2183
rect 2806 2149 2817 2183
rect 2764 2115 2817 2149
rect 2764 2081 2772 2115
rect 2806 2081 2817 2115
rect 2764 2047 2817 2081
rect 2764 2013 2772 2047
rect 2806 2013 2817 2047
rect 2764 1979 2817 2013
rect 2764 1945 2772 1979
rect 2806 1945 2817 1979
rect 2764 1911 2817 1945
rect 2764 1877 2772 1911
rect 2806 1877 2817 1911
rect 2764 1865 2817 1877
rect 2917 2795 2973 2865
rect 2917 2761 2928 2795
rect 2962 2761 2973 2795
rect 2917 2727 2973 2761
rect 2917 2693 2928 2727
rect 2962 2693 2973 2727
rect 2917 2659 2973 2693
rect 2917 2625 2928 2659
rect 2962 2625 2973 2659
rect 2917 2591 2973 2625
rect 2917 2557 2928 2591
rect 2962 2557 2973 2591
rect 2917 2523 2973 2557
rect 2917 2489 2928 2523
rect 2962 2489 2973 2523
rect 2917 2455 2973 2489
rect 2917 2421 2928 2455
rect 2962 2421 2973 2455
rect 2917 2387 2973 2421
rect 2917 2353 2928 2387
rect 2962 2353 2973 2387
rect 2917 2319 2973 2353
rect 2917 2285 2928 2319
rect 2962 2285 2973 2319
rect 2917 2251 2973 2285
rect 2917 2217 2928 2251
rect 2962 2217 2973 2251
rect 2917 2183 2973 2217
rect 2917 2149 2928 2183
rect 2962 2149 2973 2183
rect 2917 2115 2973 2149
rect 2917 2081 2928 2115
rect 2962 2081 2973 2115
rect 2917 2047 2973 2081
rect 2917 2013 2928 2047
rect 2962 2013 2973 2047
rect 2917 1979 2973 2013
rect 2917 1945 2928 1979
rect 2962 1945 2973 1979
rect 2917 1911 2973 1945
rect 2917 1877 2928 1911
rect 2962 1877 2973 1911
rect 2917 1865 2973 1877
rect 3073 2795 3126 2865
rect 3073 2761 3084 2795
rect 3118 2761 3126 2795
rect 3073 2727 3126 2761
rect 3073 2693 3084 2727
rect 3118 2693 3126 2727
rect 3073 2659 3126 2693
rect 3073 2625 3084 2659
rect 3118 2625 3126 2659
rect 3073 2591 3126 2625
rect 3073 2557 3084 2591
rect 3118 2557 3126 2591
rect 3073 2523 3126 2557
rect 3073 2489 3084 2523
rect 3118 2489 3126 2523
rect 3073 2455 3126 2489
rect 3073 2421 3084 2455
rect 3118 2421 3126 2455
rect 3073 2387 3126 2421
rect 3073 2353 3084 2387
rect 3118 2353 3126 2387
rect 3073 2319 3126 2353
rect 3073 2285 3084 2319
rect 3118 2285 3126 2319
rect 3073 2251 3126 2285
rect 3073 2217 3084 2251
rect 3118 2217 3126 2251
rect 3073 2183 3126 2217
rect 3073 2149 3084 2183
rect 3118 2149 3126 2183
rect 3073 2115 3126 2149
rect 3073 2081 3084 2115
rect 3118 2081 3126 2115
rect 3073 2047 3126 2081
rect 3073 2013 3084 2047
rect 3118 2013 3126 2047
rect 3073 1979 3126 2013
rect 3073 1945 3084 1979
rect 3118 1945 3126 1979
rect 3073 1911 3126 1945
rect 3073 1877 3084 1911
rect 3118 1877 3126 1911
rect 3073 1865 3126 1877
<< mvndiffc >>
rect 44 94 78 128
rect 44 26 78 60
rect 44 -42 78 -8
rect 44 -110 78 -76
rect 44 -178 78 -144
rect 44 -246 78 -212
rect 44 -314 78 -280
rect 44 -382 78 -348
rect 44 -450 78 -416
rect 44 -518 78 -484
rect 44 -586 78 -552
rect 44 -654 78 -620
rect 44 -722 78 -688
rect 44 -790 78 -756
rect 260 94 294 128
rect 260 26 294 60
rect 260 -42 294 -8
rect 260 -110 294 -76
rect 260 -178 294 -144
rect 260 -246 294 -212
rect 260 -314 294 -280
rect 260 -382 294 -348
rect 260 -450 294 -416
rect 260 -518 294 -484
rect 260 -586 294 -552
rect 260 -654 294 -620
rect 260 -722 294 -688
rect 260 -790 294 -756
rect 476 94 510 128
rect 476 26 510 60
rect 476 -42 510 -8
rect 476 -110 510 -76
rect 476 -178 510 -144
rect 476 -246 510 -212
rect 476 -314 510 -280
rect 476 -382 510 -348
rect 476 -450 510 -416
rect 476 -518 510 -484
rect 476 -586 510 -552
rect 476 -654 510 -620
rect 476 -722 510 -688
rect 476 -790 510 -756
rect 692 94 726 128
rect 692 26 726 60
rect 692 -42 726 -8
rect 692 -110 726 -76
rect 692 -178 726 -144
rect 692 -246 726 -212
rect 692 -314 726 -280
rect 692 -382 726 -348
rect 692 -450 726 -416
rect 692 -518 726 -484
rect 692 -586 726 -552
rect 692 -654 726 -620
rect 692 -722 726 -688
rect 692 -790 726 -756
rect 908 94 942 128
rect 908 26 942 60
rect 908 -42 942 -8
rect 908 -110 942 -76
rect 908 -178 942 -144
rect 908 -246 942 -212
rect 908 -314 942 -280
rect 908 -382 942 -348
rect 908 -450 942 -416
rect 908 -518 942 -484
rect 908 -586 942 -552
rect 908 -654 942 -620
rect 908 -722 942 -688
rect 908 -790 942 -756
rect 1124 94 1158 128
rect 1124 26 1158 60
rect 1124 -42 1158 -8
rect 1124 -110 1158 -76
rect 1124 -178 1158 -144
rect 1124 -246 1158 -212
rect 1124 -314 1158 -280
rect 1124 -382 1158 -348
rect 1124 -450 1158 -416
rect 1124 -518 1158 -484
rect 1124 -586 1158 -552
rect 1124 -654 1158 -620
rect 1124 -722 1158 -688
rect 1124 -790 1158 -756
rect 1340 94 1374 128
rect 1340 26 1374 60
rect 1340 -42 1374 -8
rect 1340 -110 1374 -76
rect 1340 -178 1374 -144
rect 1340 -246 1374 -212
rect 1340 -314 1374 -280
rect 1340 -382 1374 -348
rect 1340 -450 1374 -416
rect 1340 -518 1374 -484
rect 1340 -586 1374 -552
rect 1340 -654 1374 -620
rect 1340 -722 1374 -688
rect 1340 -790 1374 -756
rect 1556 94 1590 128
rect 1556 26 1590 60
rect 1556 -42 1590 -8
rect 1556 -110 1590 -76
rect 1556 -178 1590 -144
rect 1556 -246 1590 -212
rect 1556 -314 1590 -280
rect 1556 -382 1590 -348
rect 1556 -450 1590 -416
rect 1556 -518 1590 -484
rect 1556 -586 1590 -552
rect 1556 -654 1590 -620
rect 1556 -722 1590 -688
rect 1556 -790 1590 -756
rect 1772 94 1806 128
rect 1772 26 1806 60
rect 1772 -42 1806 -8
rect 1772 -110 1806 -76
rect 1772 -178 1806 -144
rect 1772 -246 1806 -212
rect 1772 -314 1806 -280
rect 1772 -382 1806 -348
rect 1772 -450 1806 -416
rect 1772 -518 1806 -484
rect 1772 -586 1806 -552
rect 1772 -654 1806 -620
rect 1772 -722 1806 -688
rect 1772 -790 1806 -756
rect 1988 94 2022 128
rect 1988 26 2022 60
rect 1988 -42 2022 -8
rect 1988 -110 2022 -76
rect 1988 -178 2022 -144
rect 1988 -246 2022 -212
rect 1988 -314 2022 -280
rect 1988 -382 2022 -348
rect 1988 -450 2022 -416
rect 1988 -518 2022 -484
rect 1988 -586 2022 -552
rect 1988 -654 2022 -620
rect 1988 -722 2022 -688
rect 1988 -790 2022 -756
rect 2204 94 2238 128
rect 2204 26 2238 60
rect 2204 -42 2238 -8
rect 2204 -110 2238 -76
rect 2204 -178 2238 -144
rect 2204 -246 2238 -212
rect 2204 -314 2238 -280
rect 2204 -382 2238 -348
rect 2204 -450 2238 -416
rect 2204 -518 2238 -484
rect 2204 -586 2238 -552
rect 2204 -654 2238 -620
rect 2204 -722 2238 -688
rect 2204 -790 2238 -756
rect 2420 94 2454 128
rect 2420 26 2454 60
rect 2420 -42 2454 -8
rect 2420 -110 2454 -76
rect 2420 -178 2454 -144
rect 2420 -246 2454 -212
rect 2420 -314 2454 -280
rect 2420 -382 2454 -348
rect 2420 -450 2454 -416
rect 2420 -518 2454 -484
rect 2420 -586 2454 -552
rect 2420 -654 2454 -620
rect 2420 -722 2454 -688
rect 2420 -790 2454 -756
rect 2636 94 2670 128
rect 2636 26 2670 60
rect 2636 -42 2670 -8
rect 2636 -110 2670 -76
rect 2636 -178 2670 -144
rect 2636 -246 2670 -212
rect 2636 -314 2670 -280
rect 2636 -382 2670 -348
rect 2636 -450 2670 -416
rect 2636 -518 2670 -484
rect 2636 -586 2670 -552
rect 2636 -654 2670 -620
rect 2636 -722 2670 -688
rect 2636 -790 2670 -756
rect 2852 94 2886 128
rect 2852 26 2886 60
rect 2852 -42 2886 -8
rect 2852 -110 2886 -76
rect 2852 -178 2886 -144
rect 2852 -246 2886 -212
rect 2852 -314 2886 -280
rect 2852 -382 2886 -348
rect 2852 -450 2886 -416
rect 2852 -518 2886 -484
rect 2852 -586 2886 -552
rect 2852 -654 2886 -620
rect 2852 -722 2886 -688
rect 2852 -790 2886 -756
rect 3068 94 3102 128
rect 3068 26 3102 60
rect 3068 -42 3102 -8
rect 3068 -110 3102 -76
rect 3068 -178 3102 -144
rect 3068 -246 3102 -212
rect 3068 -314 3102 -280
rect 3068 -382 3102 -348
rect 3068 -450 3102 -416
rect 3068 -518 3102 -484
rect 3068 -586 3102 -552
rect 3068 -654 3102 -620
rect 3068 -722 3102 -688
rect 3068 -790 3102 -756
rect 3284 94 3318 128
rect 3284 26 3318 60
rect 3284 -42 3318 -8
rect 3284 -110 3318 -76
rect 3284 -178 3318 -144
rect 3284 -246 3318 -212
rect 3284 -314 3318 -280
rect 3284 -382 3318 -348
rect 3284 -450 3318 -416
rect 3284 -518 3318 -484
rect 3284 -586 3318 -552
rect 3284 -654 3318 -620
rect 3284 -722 3318 -688
rect 3284 -790 3318 -756
rect 3394 94 3428 128
rect 3394 26 3428 60
rect 3394 -42 3428 -8
rect 3394 -110 3428 -76
rect 3394 -178 3428 -144
rect 3394 -246 3428 -212
rect 3394 -314 3428 -280
rect 3394 -382 3428 -348
rect 3394 -450 3428 -416
rect 3394 -518 3428 -484
rect 3394 -586 3428 -552
rect 3394 -654 3428 -620
rect 3394 -722 3428 -688
rect 3394 -790 3428 -756
rect 3610 94 3644 128
rect 3610 26 3644 60
rect 3610 -42 3644 -8
rect 3610 -110 3644 -76
rect 3610 -178 3644 -144
rect 3610 -246 3644 -212
rect 3610 -314 3644 -280
rect 3610 -382 3644 -348
rect 3610 -450 3644 -416
rect 3610 -518 3644 -484
rect 3610 -586 3644 -552
rect 3610 -654 3644 -620
rect 3610 -722 3644 -688
rect 3610 -790 3644 -756
rect 3720 94 3754 128
rect 3720 26 3754 60
rect 3720 -42 3754 -8
rect 3720 -110 3754 -76
rect 3720 -178 3754 -144
rect 3720 -246 3754 -212
rect 3720 -314 3754 -280
rect 3720 -382 3754 -348
rect 3720 -450 3754 -416
rect 3720 -518 3754 -484
rect 3720 -586 3754 -552
rect 3720 -654 3754 -620
rect 3720 -722 3754 -688
rect 3720 -790 3754 -756
rect 3936 94 3970 128
rect 3936 26 3970 60
rect 3936 -42 3970 -8
rect 3936 -110 3970 -76
rect 3936 -178 3970 -144
rect 3936 -246 3970 -212
rect 3936 -314 3970 -280
rect 3936 -382 3970 -348
rect 3936 -450 3970 -416
rect 3936 -518 3970 -484
rect 3936 -586 3970 -552
rect 3936 -654 3970 -620
rect 3936 -722 3970 -688
rect 3936 -790 3970 -756
rect 4046 94 4080 128
rect 4046 26 4080 60
rect 4046 -42 4080 -8
rect 4046 -110 4080 -76
rect 4046 -178 4080 -144
rect 4046 -246 4080 -212
rect 4046 -314 4080 -280
rect 4046 -382 4080 -348
rect 4046 -450 4080 -416
rect 4046 -518 4080 -484
rect 4046 -586 4080 -552
rect 4046 -654 4080 -620
rect 4046 -722 4080 -688
rect 4046 -790 4080 -756
rect 4262 94 4296 128
rect 4262 26 4296 60
rect 4372 167 4406 201
rect 4372 99 4406 133
rect 4372 31 4406 65
rect 4588 167 4622 201
rect 4588 99 4622 133
rect 4588 31 4622 65
rect 4804 167 4838 201
rect 4804 99 4838 133
rect 4804 31 4838 65
rect 5020 167 5054 201
rect 5020 99 5054 133
rect 5020 31 5054 65
rect 5236 167 5270 201
rect 5236 99 5270 133
rect 5236 31 5270 65
rect 5362 94 5396 128
rect 5362 26 5396 60
rect 4262 -42 4296 -8
rect 4262 -110 4296 -76
rect 5362 -42 5396 -8
rect 4262 -178 4296 -144
rect 5362 -110 5396 -76
rect 5362 -178 5396 -144
rect 4262 -246 4296 -212
rect 4262 -314 4296 -280
rect 4262 -382 4296 -348
rect 4262 -450 4296 -416
rect 4262 -518 4296 -484
rect 4262 -586 4296 -552
rect 4262 -654 4296 -620
rect 4262 -722 4296 -688
rect 4262 -790 4296 -756
rect 4372 -314 4406 -280
rect 4372 -382 4406 -348
rect 4372 -450 4406 -416
rect 4372 -518 4406 -484
rect 4372 -586 4406 -552
rect 4372 -654 4406 -620
rect 4372 -722 4406 -688
rect 4372 -790 4406 -756
rect 4628 -314 4662 -280
rect 4628 -382 4662 -348
rect 4628 -450 4662 -416
rect 4628 -518 4662 -484
rect 4628 -586 4662 -552
rect 4628 -654 4662 -620
rect 4628 -722 4662 -688
rect 4628 -790 4662 -756
rect 4784 -314 4818 -280
rect 4784 -382 4818 -348
rect 4784 -450 4818 -416
rect 4784 -518 4818 -484
rect 4784 -586 4818 -552
rect 4784 -654 4818 -620
rect 4784 -722 4818 -688
rect 4784 -790 4818 -756
rect 4940 -314 4974 -280
rect 4940 -382 4974 -348
rect 4940 -450 4974 -416
rect 4940 -518 4974 -484
rect 4940 -586 4974 -552
rect 4940 -654 4974 -620
rect 4940 -722 4974 -688
rect 4940 -790 4974 -756
rect 5096 -314 5130 -280
rect 5096 -382 5130 -348
rect 5096 -450 5130 -416
rect 5096 -518 5130 -484
rect 5096 -586 5130 -552
rect 5096 -654 5130 -620
rect 5096 -722 5130 -688
rect 5096 -790 5130 -756
rect 5252 -314 5286 -280
rect 5252 -382 5286 -348
rect 5252 -450 5286 -416
rect 5252 -518 5286 -484
rect 5252 -586 5286 -552
rect 5252 -654 5286 -620
rect 5252 -722 5286 -688
rect 5252 -790 5286 -756
rect 5362 -246 5396 -212
rect 5362 -314 5396 -280
rect 5362 -382 5396 -348
rect 5362 -450 5396 -416
rect 5362 -518 5396 -484
rect 5362 -586 5396 -552
rect 5362 -654 5396 -620
rect 5362 -722 5396 -688
rect 5362 -790 5396 -756
rect 5518 94 5552 128
rect 5518 26 5552 60
rect 5518 -42 5552 -8
rect 5518 -110 5552 -76
rect 5518 -178 5552 -144
rect 5518 -246 5552 -212
rect 5518 -314 5552 -280
rect 5518 -382 5552 -348
rect 5518 -450 5552 -416
rect 5518 -518 5552 -484
rect 5518 -586 5552 -552
rect 5518 -654 5552 -620
rect 5518 -722 5552 -688
rect 5518 -790 5552 -756
rect 5674 94 5708 128
rect 5674 26 5708 60
rect 5674 -42 5708 -8
rect 5674 -110 5708 -76
rect 5674 -178 5708 -144
rect 5674 -246 5708 -212
rect 5674 -314 5708 -280
rect 5674 -382 5708 -348
rect 5674 -450 5708 -416
rect 5674 -518 5708 -484
rect 5674 -586 5708 -552
rect 5674 -654 5708 -620
rect 5674 -722 5708 -688
rect 5674 -790 5708 -756
<< mvpdiffc >>
rect 74 2761 108 2795
rect 74 2693 108 2727
rect 74 2625 108 2659
rect 74 2557 108 2591
rect 74 2489 108 2523
rect 74 2421 108 2455
rect 74 2353 108 2387
rect 74 2285 108 2319
rect 74 2217 108 2251
rect 74 2149 108 2183
rect 74 2081 108 2115
rect 74 2013 108 2047
rect 74 1945 108 1979
rect 74 1877 108 1911
rect 230 2761 264 2795
rect 230 2693 264 2727
rect 230 2625 264 2659
rect 230 2557 264 2591
rect 230 2489 264 2523
rect 230 2421 264 2455
rect 230 2353 264 2387
rect 230 2285 264 2319
rect 230 2217 264 2251
rect 230 2149 264 2183
rect 230 2081 264 2115
rect 230 2013 264 2047
rect 230 1945 264 1979
rect 230 1877 264 1911
rect 386 2761 420 2795
rect 386 2693 420 2727
rect 386 2625 420 2659
rect 386 2557 420 2591
rect 386 2489 420 2523
rect 386 2421 420 2455
rect 386 2353 420 2387
rect 386 2285 420 2319
rect 386 2217 420 2251
rect 386 2149 420 2183
rect 386 2081 420 2115
rect 386 2013 420 2047
rect 386 1945 420 1979
rect 386 1877 420 1911
rect 496 2761 530 2795
rect 496 2693 530 2727
rect 496 2625 530 2659
rect 496 2557 530 2591
rect 496 2489 530 2523
rect 496 2421 530 2455
rect 496 2353 530 2387
rect 496 2285 530 2319
rect 496 2217 530 2251
rect 496 2149 530 2183
rect 496 2081 530 2115
rect 496 2013 530 2047
rect 496 1945 530 1979
rect 496 1877 530 1911
rect 712 2761 746 2795
rect 712 2693 746 2727
rect 712 2625 746 2659
rect 712 2557 746 2591
rect 712 2489 746 2523
rect 712 2421 746 2455
rect 712 2353 746 2387
rect 712 2285 746 2319
rect 712 2217 746 2251
rect 712 2149 746 2183
rect 712 2081 746 2115
rect 712 2013 746 2047
rect 712 1945 746 1979
rect 712 1877 746 1911
rect 928 2761 962 2795
rect 928 2693 962 2727
rect 928 2625 962 2659
rect 928 2557 962 2591
rect 928 2489 962 2523
rect 928 2421 962 2455
rect 928 2353 962 2387
rect 928 2285 962 2319
rect 928 2217 962 2251
rect 928 2149 962 2183
rect 928 2081 962 2115
rect 928 2013 962 2047
rect 928 1945 962 1979
rect 928 1877 962 1911
rect 1084 2761 1118 2795
rect 1084 2693 1118 2727
rect 1084 2625 1118 2659
rect 1084 2557 1118 2591
rect 1084 2489 1118 2523
rect 1084 2421 1118 2455
rect 1084 2353 1118 2387
rect 1084 2285 1118 2319
rect 1084 2217 1118 2251
rect 1084 2149 1118 2183
rect 1084 2081 1118 2115
rect 1084 2013 1118 2047
rect 1084 1945 1118 1979
rect 1084 1877 1118 1911
rect 1240 2761 1274 2795
rect 1240 2693 1274 2727
rect 1240 2625 1274 2659
rect 1240 2557 1274 2591
rect 1240 2489 1274 2523
rect 1240 2421 1274 2455
rect 1240 2353 1274 2387
rect 1240 2285 1274 2319
rect 1240 2217 1274 2251
rect 1240 2149 1274 2183
rect 1240 2081 1274 2115
rect 1240 2013 1274 2047
rect 1240 1945 1274 1979
rect 1240 1877 1274 1911
rect 1400 2761 1434 2795
rect 1400 2693 1434 2727
rect 1400 2625 1434 2659
rect 1400 2557 1434 2591
rect 1400 2489 1434 2523
rect 1400 2421 1434 2455
rect 1400 2353 1434 2387
rect 1400 2285 1434 2319
rect 1400 2217 1434 2251
rect 1400 2149 1434 2183
rect 1400 2081 1434 2115
rect 1400 2013 1434 2047
rect 1400 1945 1434 1979
rect 1400 1877 1434 1911
rect 1616 2761 1650 2795
rect 1616 2693 1650 2727
rect 1616 2625 1650 2659
rect 1616 2557 1650 2591
rect 1616 2489 1650 2523
rect 1616 2421 1650 2455
rect 1616 2353 1650 2387
rect 1616 2285 1650 2319
rect 1616 2217 1650 2251
rect 1616 2149 1650 2183
rect 1616 2081 1650 2115
rect 1616 2013 1650 2047
rect 1616 1945 1650 1979
rect 1616 1877 1650 1911
rect 1772 2761 1806 2795
rect 1772 2693 1806 2727
rect 1772 2625 1806 2659
rect 1772 2557 1806 2591
rect 1772 2489 1806 2523
rect 1772 2421 1806 2455
rect 1772 2353 1806 2387
rect 1772 2285 1806 2319
rect 1772 2217 1806 2251
rect 1772 2149 1806 2183
rect 1772 2081 1806 2115
rect 1772 2013 1806 2047
rect 1772 1945 1806 1979
rect 1772 1877 1806 1911
rect 1928 2761 1962 2795
rect 1928 2693 1962 2727
rect 1928 2625 1962 2659
rect 1928 2557 1962 2591
rect 1928 2489 1962 2523
rect 1928 2421 1962 2455
rect 1928 2353 1962 2387
rect 1928 2285 1962 2319
rect 1928 2217 1962 2251
rect 1928 2149 1962 2183
rect 1928 2081 1962 2115
rect 1928 2013 1962 2047
rect 1928 1945 1962 1979
rect 1928 1877 1962 1911
rect 2084 2761 2118 2795
rect 2084 2693 2118 2727
rect 2084 2625 2118 2659
rect 2084 2557 2118 2591
rect 2084 2489 2118 2523
rect 2084 2421 2118 2455
rect 2084 2353 2118 2387
rect 2084 2285 2118 2319
rect 2084 2217 2118 2251
rect 2084 2149 2118 2183
rect 2084 2081 2118 2115
rect 2084 2013 2118 2047
rect 2084 1945 2118 1979
rect 2084 1877 2118 1911
rect 2240 2761 2274 2795
rect 2240 2693 2274 2727
rect 2240 2625 2274 2659
rect 2240 2557 2274 2591
rect 2240 2489 2274 2523
rect 2240 2421 2274 2455
rect 2240 2353 2274 2387
rect 2240 2285 2274 2319
rect 2240 2217 2274 2251
rect 2240 2149 2274 2183
rect 2240 2081 2274 2115
rect 2240 2013 2274 2047
rect 2240 1945 2274 1979
rect 2240 1877 2274 1911
rect 2396 2761 2430 2795
rect 2396 2693 2430 2727
rect 2396 2625 2430 2659
rect 2396 2557 2430 2591
rect 2396 2489 2430 2523
rect 2772 2761 2806 2795
rect 2772 2693 2806 2727
rect 2772 2625 2806 2659
rect 2772 2557 2806 2591
rect 2772 2489 2806 2523
rect 2396 2421 2430 2455
rect 2396 2353 2430 2387
rect 2396 2285 2430 2319
rect 2396 2217 2430 2251
rect 2396 2149 2430 2183
rect 2396 2081 2430 2115
rect 2396 2013 2430 2047
rect 2396 1945 2430 1979
rect 2396 1877 2430 1911
rect 2506 2353 2540 2387
rect 2506 2285 2540 2319
rect 2506 2217 2540 2251
rect 2506 2149 2540 2183
rect 2506 2081 2540 2115
rect 2506 2013 2540 2047
rect 2506 1945 2540 1979
rect 2506 1877 2540 1911
rect 2662 2353 2696 2387
rect 2662 2285 2696 2319
rect 2662 2217 2696 2251
rect 2662 2149 2696 2183
rect 2662 2081 2696 2115
rect 2662 2013 2696 2047
rect 2662 1945 2696 1979
rect 2662 1877 2696 1911
rect 2772 2421 2806 2455
rect 2772 2353 2806 2387
rect 2772 2285 2806 2319
rect 2772 2217 2806 2251
rect 2772 2149 2806 2183
rect 2772 2081 2806 2115
rect 2772 2013 2806 2047
rect 2772 1945 2806 1979
rect 2772 1877 2806 1911
rect 2928 2761 2962 2795
rect 2928 2693 2962 2727
rect 2928 2625 2962 2659
rect 2928 2557 2962 2591
rect 2928 2489 2962 2523
rect 2928 2421 2962 2455
rect 2928 2353 2962 2387
rect 2928 2285 2962 2319
rect 2928 2217 2962 2251
rect 2928 2149 2962 2183
rect 2928 2081 2962 2115
rect 2928 2013 2962 2047
rect 2928 1945 2962 1979
rect 2928 1877 2962 1911
rect 3084 2761 3118 2795
rect 3084 2693 3118 2727
rect 3084 2625 3118 2659
rect 3084 2557 3118 2591
rect 3084 2489 3118 2523
rect 3084 2421 3118 2455
rect 3084 2353 3118 2387
rect 3084 2285 3118 2319
rect 3084 2217 3118 2251
rect 3084 2149 3118 2183
rect 3084 2081 3118 2115
rect 3084 2013 3118 2047
rect 3084 1945 3118 1979
rect 3084 1877 3118 1911
<< mvpsubdiff >>
rect 67 -912 91 -878
rect 125 -912 160 -878
rect 194 -912 229 -878
rect 263 -912 298 -878
rect 332 -912 367 -878
rect 401 -912 436 -878
rect 470 -912 505 -878
rect 539 -912 574 -878
rect 608 -912 643 -878
rect 677 -912 712 -878
rect 746 -912 781 -878
rect 815 -912 850 -878
rect 884 -912 919 -878
rect 953 -912 988 -878
rect 1022 -912 1057 -878
rect 1091 -912 1126 -878
rect 1160 -912 1195 -878
rect 1229 -912 1264 -878
rect 1298 -912 1333 -878
rect 1367 -912 1402 -878
rect 1436 -912 1471 -878
rect 1505 -912 1540 -878
rect 1574 -912 1609 -878
rect 1643 -912 1678 -878
rect 1712 -912 1747 -878
rect 1781 -912 1816 -878
rect 1850 -912 1885 -878
rect 1919 -912 1954 -878
rect 1988 -912 2023 -878
rect 2057 -912 2092 -878
rect 2126 -912 2161 -878
rect 2195 -912 2230 -878
rect 2264 -912 2299 -878
rect 2333 -912 2368 -878
rect 2402 -912 2437 -878
rect 2471 -912 2505 -878
rect 2539 -912 2573 -878
rect 2607 -912 2641 -878
rect 2675 -912 2709 -878
rect 2743 -912 2777 -878
rect 2811 -912 2845 -878
rect 2879 -912 2913 -878
rect 2947 -912 2981 -878
rect 3015 -912 3049 -878
rect 3083 -912 3117 -878
rect 3151 -912 3185 -878
rect 3219 -912 3253 -878
rect 3287 -912 3321 -878
rect 3355 -912 3389 -878
rect 3423 -912 3457 -878
rect 3491 -912 3525 -878
rect 3559 -912 3593 -878
rect 3627 -912 3661 -878
rect 3695 -912 3729 -878
rect 3763 -912 3797 -878
rect 3831 -912 3865 -878
rect 3899 -912 3933 -878
rect 3967 -912 4001 -878
rect 4035 -912 4069 -878
rect 4103 -912 4137 -878
rect 4171 -912 4205 -878
rect 4239 -912 4273 -878
rect 4307 -912 4341 -878
rect 4375 -912 4409 -878
rect 4443 -912 4477 -878
rect 4511 -912 4545 -878
rect 4579 -912 4613 -878
rect 4647 -912 4681 -878
rect 4715 -912 4749 -878
rect 4783 -912 4817 -878
rect 4851 -912 4885 -878
rect 4919 -912 4953 -878
rect 4987 -912 5021 -878
rect 5055 -912 5089 -878
rect 5123 -912 5157 -878
rect 5191 -912 5225 -878
rect 5259 -912 5293 -878
rect 5327 -912 5361 -878
rect 5395 -912 5429 -878
rect 5463 -912 5497 -878
rect 5531 -912 5565 -878
rect 5599 -912 5633 -878
rect 5667 -912 5691 -878
<< mvnsubdiff >>
rect 67 2947 101 2981
rect 135 2947 169 2981
rect 203 2947 237 2981
rect 271 2947 305 2981
rect 339 2947 373 2981
rect 407 2947 441 2981
rect 475 2947 509 2981
rect 543 2947 577 2981
rect 611 2947 645 2981
rect 679 2947 713 2981
rect 747 2947 781 2981
rect 815 2947 849 2981
rect 883 2947 917 2981
rect 951 2947 985 2981
rect 1019 2947 1053 2981
rect 1087 2947 1121 2981
rect 1155 2947 1189 2981
rect 1223 2947 1257 2981
rect 1291 2947 1325 2981
rect 1359 2947 1393 2981
rect 1427 2947 1461 2981
rect 1495 2947 1529 2981
rect 1563 2947 1597 2981
rect 1631 2947 1665 2981
rect 1699 2947 1733 2981
rect 1767 2947 1801 2981
rect 1835 2947 1869 2981
rect 1903 2947 1937 2981
rect 1971 2947 2005 2981
rect 2039 2947 2073 2981
rect 2107 2947 2141 2981
rect 2175 2947 2209 2981
rect 2243 2947 2277 2981
rect 2311 2947 2345 2981
rect 2379 2947 2413 2981
rect 2447 2947 2481 2981
rect 2515 2947 2549 2981
rect 2583 2947 2617 2981
rect 2651 2947 2685 2981
rect 2719 2947 2753 2981
rect 2787 2947 2821 2981
rect 2855 2947 2889 2981
rect 2923 2947 2957 2981
rect 2991 2947 3025 2981
rect 3059 2947 3093 2981
rect 3127 2947 3161 2981
rect 3195 2947 3229 2981
rect 3263 2947 3297 2981
rect 3331 2947 3365 2981
rect 3399 2947 3433 2981
rect 3467 2947 3501 2981
rect 3535 2947 3569 2981
rect 3603 2947 3637 2981
rect 3671 2947 3705 2981
rect 3739 2947 3773 2981
rect 3807 2947 3841 2981
rect 3875 2947 3976 2981
<< mvpsubdiffcont >>
rect 91 -912 125 -878
rect 160 -912 194 -878
rect 229 -912 263 -878
rect 298 -912 332 -878
rect 367 -912 401 -878
rect 436 -912 470 -878
rect 505 -912 539 -878
rect 574 -912 608 -878
rect 643 -912 677 -878
rect 712 -912 746 -878
rect 781 -912 815 -878
rect 850 -912 884 -878
rect 919 -912 953 -878
rect 988 -912 1022 -878
rect 1057 -912 1091 -878
rect 1126 -912 1160 -878
rect 1195 -912 1229 -878
rect 1264 -912 1298 -878
rect 1333 -912 1367 -878
rect 1402 -912 1436 -878
rect 1471 -912 1505 -878
rect 1540 -912 1574 -878
rect 1609 -912 1643 -878
rect 1678 -912 1712 -878
rect 1747 -912 1781 -878
rect 1816 -912 1850 -878
rect 1885 -912 1919 -878
rect 1954 -912 1988 -878
rect 2023 -912 2057 -878
rect 2092 -912 2126 -878
rect 2161 -912 2195 -878
rect 2230 -912 2264 -878
rect 2299 -912 2333 -878
rect 2368 -912 2402 -878
rect 2437 -912 2471 -878
rect 2505 -912 2539 -878
rect 2573 -912 2607 -878
rect 2641 -912 2675 -878
rect 2709 -912 2743 -878
rect 2777 -912 2811 -878
rect 2845 -912 2879 -878
rect 2913 -912 2947 -878
rect 2981 -912 3015 -878
rect 3049 -912 3083 -878
rect 3117 -912 3151 -878
rect 3185 -912 3219 -878
rect 3253 -912 3287 -878
rect 3321 -912 3355 -878
rect 3389 -912 3423 -878
rect 3457 -912 3491 -878
rect 3525 -912 3559 -878
rect 3593 -912 3627 -878
rect 3661 -912 3695 -878
rect 3729 -912 3763 -878
rect 3797 -912 3831 -878
rect 3865 -912 3899 -878
rect 3933 -912 3967 -878
rect 4001 -912 4035 -878
rect 4069 -912 4103 -878
rect 4137 -912 4171 -878
rect 4205 -912 4239 -878
rect 4273 -912 4307 -878
rect 4341 -912 4375 -878
rect 4409 -912 4443 -878
rect 4477 -912 4511 -878
rect 4545 -912 4579 -878
rect 4613 -912 4647 -878
rect 4681 -912 4715 -878
rect 4749 -912 4783 -878
rect 4817 -912 4851 -878
rect 4885 -912 4919 -878
rect 4953 -912 4987 -878
rect 5021 -912 5055 -878
rect 5089 -912 5123 -878
rect 5157 -912 5191 -878
rect 5225 -912 5259 -878
rect 5293 -912 5327 -878
rect 5361 -912 5395 -878
rect 5429 -912 5463 -878
rect 5497 -912 5531 -878
rect 5565 -912 5599 -878
rect 5633 -912 5667 -878
<< mvnsubdiffcont >>
rect 101 2947 135 2981
rect 169 2947 203 2981
rect 237 2947 271 2981
rect 305 2947 339 2981
rect 373 2947 407 2981
rect 441 2947 475 2981
rect 509 2947 543 2981
rect 577 2947 611 2981
rect 645 2947 679 2981
rect 713 2947 747 2981
rect 781 2947 815 2981
rect 849 2947 883 2981
rect 917 2947 951 2981
rect 985 2947 1019 2981
rect 1053 2947 1087 2981
rect 1121 2947 1155 2981
rect 1189 2947 1223 2981
rect 1257 2947 1291 2981
rect 1325 2947 1359 2981
rect 1393 2947 1427 2981
rect 1461 2947 1495 2981
rect 1529 2947 1563 2981
rect 1597 2947 1631 2981
rect 1665 2947 1699 2981
rect 1733 2947 1767 2981
rect 1801 2947 1835 2981
rect 1869 2947 1903 2981
rect 1937 2947 1971 2981
rect 2005 2947 2039 2981
rect 2073 2947 2107 2981
rect 2141 2947 2175 2981
rect 2209 2947 2243 2981
rect 2277 2947 2311 2981
rect 2345 2947 2379 2981
rect 2413 2947 2447 2981
rect 2481 2947 2515 2981
rect 2549 2947 2583 2981
rect 2617 2947 2651 2981
rect 2685 2947 2719 2981
rect 2753 2947 2787 2981
rect 2821 2947 2855 2981
rect 2889 2947 2923 2981
rect 2957 2947 2991 2981
rect 3025 2947 3059 2981
rect 3093 2947 3127 2981
rect 3161 2947 3195 2981
rect 3229 2947 3263 2981
rect 3297 2947 3331 2981
rect 3365 2947 3399 2981
rect 3433 2947 3467 2981
rect 3501 2947 3535 2981
rect 3569 2947 3603 2981
rect 3637 2947 3671 2981
rect 3705 2947 3739 2981
rect 3773 2947 3807 2981
rect 3841 2947 3875 2981
<< poly >>
rect 119 2865 219 2897
rect 275 2865 375 2897
rect 541 2865 701 2897
rect 757 2865 917 2897
rect 973 2865 1073 2897
rect 1129 2865 1229 2897
rect 1445 2865 1605 2897
rect 1661 2865 1761 2897
rect 1817 2865 1917 2897
rect 1973 2865 2073 2897
rect 2129 2865 2229 2897
rect 2285 2865 2385 2897
rect 2817 2865 2917 2897
rect 2973 2865 3073 2897
rect 2551 2465 2651 2497
rect 119 1833 219 1865
rect 275 1833 375 1865
rect 119 1817 375 1833
rect 119 1783 135 1817
rect 169 1783 230 1817
rect 264 1783 325 1817
rect 359 1783 375 1817
rect 119 1767 375 1783
rect 541 1817 701 1865
rect 541 1783 557 1817
rect 591 1783 651 1817
rect 685 1783 701 1817
rect 541 1767 701 1783
rect 757 1817 917 1865
rect 757 1783 773 1817
rect 807 1783 867 1817
rect 901 1783 917 1817
rect 757 1767 917 1783
rect 973 1833 1073 1865
rect 1129 1833 1229 1865
rect 1445 1833 1605 1865
rect 973 1817 1229 1833
rect 973 1783 989 1817
rect 1023 1783 1084 1817
rect 1118 1783 1179 1817
rect 1213 1783 1229 1817
rect 973 1767 1229 1783
rect 1471 1817 1605 1833
rect 1471 1783 1487 1817
rect 1521 1783 1555 1817
rect 1589 1783 1605 1817
rect 1471 1767 1605 1783
rect 1661 1833 1761 1865
rect 1817 1833 1917 1865
rect 1661 1817 1917 1833
rect 1661 1783 1677 1817
rect 1711 1783 1772 1817
rect 1806 1783 1867 1817
rect 1901 1783 1917 1817
rect 1661 1767 1917 1783
rect 1973 1833 2073 1865
rect 2129 1833 2229 1865
rect 1973 1817 2229 1833
rect 1973 1783 1989 1817
rect 2023 1783 2084 1817
rect 2118 1783 2179 1817
rect 2213 1783 2229 1817
rect 1973 1767 2229 1783
rect 2285 1833 2385 1865
rect 2551 1833 2651 1865
rect 2817 1833 2917 1865
rect 2285 1817 2419 1833
rect 2285 1783 2301 1817
rect 2335 1783 2369 1817
rect 2403 1783 2419 1817
rect 2285 1767 2419 1783
rect 2517 1817 2651 1833
rect 2517 1783 2533 1817
rect 2567 1783 2601 1817
rect 2635 1783 2651 1817
rect 2517 1767 2651 1783
rect 2783 1817 2917 1833
rect 2783 1783 2799 1817
rect 2833 1783 2867 1817
rect 2901 1783 2917 1817
rect 2783 1767 2917 1783
rect 2973 1833 3073 1865
rect 2973 1817 3107 1833
rect 2973 1783 2989 1817
rect 3023 1783 3057 1817
rect 3091 1783 3107 1817
rect 2973 1767 3107 1783
rect 89 280 1113 296
rect 89 246 105 280
rect 139 246 174 280
rect 208 246 243 280
rect 277 246 312 280
rect 346 246 381 280
rect 415 246 450 280
rect 484 246 519 280
rect 553 246 587 280
rect 621 246 655 280
rect 689 246 723 280
rect 757 246 791 280
rect 825 246 859 280
rect 893 246 927 280
rect 961 246 995 280
rect 1029 246 1063 280
rect 1097 246 1113 280
rect 89 230 1113 246
rect 89 198 249 230
rect 305 198 465 230
rect 521 198 681 230
rect 737 198 897 230
rect 953 198 1113 230
rect 1169 280 1329 296
rect 1169 246 1185 280
rect 1219 246 1279 280
rect 1313 246 1329 280
rect 1169 198 1329 246
rect 1385 280 2409 296
rect 1385 246 1401 280
rect 1435 246 1470 280
rect 1504 246 1539 280
rect 1573 246 1608 280
rect 1642 246 1677 280
rect 1711 246 1746 280
rect 1780 246 1815 280
rect 1849 246 1883 280
rect 1917 246 1951 280
rect 1985 246 2019 280
rect 2053 246 2087 280
rect 2121 246 2155 280
rect 2189 246 2223 280
rect 2257 246 2291 280
rect 2325 246 2359 280
rect 2393 246 2409 280
rect 1385 230 2409 246
rect 1385 198 1545 230
rect 1601 198 1761 230
rect 1817 198 1977 230
rect 2033 198 2193 230
rect 2249 198 2409 230
rect 2465 280 3273 296
rect 2465 246 2481 280
rect 2515 246 2556 280
rect 2590 246 2631 280
rect 2665 246 2705 280
rect 2739 246 2779 280
rect 2813 246 2853 280
rect 2887 246 2927 280
rect 2961 246 3001 280
rect 3035 246 3075 280
rect 3109 246 3149 280
rect 3183 246 3223 280
rect 3257 246 3273 280
rect 2465 230 3273 246
rect 2465 198 2625 230
rect 2681 198 2841 230
rect 2897 198 3057 230
rect 3113 198 3273 230
rect 3439 280 3599 296
rect 3439 246 3455 280
rect 3489 246 3549 280
rect 3583 246 3599 280
rect 3439 198 3599 246
rect 3765 280 3925 296
rect 3765 246 3781 280
rect 3815 246 3875 280
rect 3909 246 3925 280
rect 3765 198 3925 246
rect 4091 280 4251 296
rect 4091 246 4107 280
rect 4141 246 4201 280
rect 4235 246 4251 280
rect 4091 198 4251 246
rect 4417 292 5225 308
rect 4417 258 4433 292
rect 4467 258 4508 292
rect 4542 258 4583 292
rect 4617 258 4657 292
rect 4691 258 4731 292
rect 4765 258 4805 292
rect 4839 258 4879 292
rect 4913 258 4953 292
rect 4987 258 5027 292
rect 5061 258 5101 292
rect 5135 258 5175 292
rect 5209 258 5225 292
rect 4417 242 5225 258
rect 4417 213 4577 242
rect 4633 213 4793 242
rect 4849 213 5009 242
rect 5065 213 5225 242
rect 5373 280 5507 296
rect 5373 246 5389 280
rect 5423 246 5457 280
rect 5491 246 5507 280
rect 5373 230 5507 246
rect 5407 198 5507 230
rect 5563 280 5697 296
rect 5563 246 5579 280
rect 5613 246 5647 280
rect 5681 246 5697 280
rect 5563 230 5697 246
rect 5563 198 5663 230
rect 4417 -19 4577 13
rect 4633 -19 4793 13
rect 4849 -19 5009 13
rect 5065 -19 5225 13
rect 4417 -120 4617 -104
rect 4417 -154 4433 -120
rect 4467 -154 4567 -120
rect 4601 -154 4617 -120
rect 4417 -202 4617 -154
rect 4673 -120 4929 -104
rect 4673 -154 4689 -120
rect 4723 -154 4784 -120
rect 4818 -154 4879 -120
rect 4913 -154 4929 -120
rect 4673 -170 4929 -154
rect 4673 -202 4773 -170
rect 4829 -202 4929 -170
rect 4985 -120 5241 -104
rect 4985 -154 5001 -120
rect 5035 -154 5096 -120
rect 5130 -154 5191 -120
rect 5225 -154 5241 -120
rect 4985 -170 5241 -154
rect 4985 -202 5085 -170
rect 5141 -202 5241 -170
rect 89 -834 249 -802
rect 305 -834 465 -802
rect 521 -834 681 -802
rect 737 -834 897 -802
rect 953 -834 1113 -802
rect 1169 -834 1329 -802
rect 1385 -834 1545 -802
rect 1601 -834 1761 -802
rect 1817 -834 1977 -802
rect 2033 -834 2193 -802
rect 2249 -834 2409 -802
rect 2465 -834 2625 -802
rect 2681 -834 2841 -802
rect 2897 -834 3057 -802
rect 3113 -834 3273 -802
rect 3439 -834 3599 -802
rect 3765 -834 3925 -802
rect 4091 -834 4251 -802
rect 4417 -834 4617 -802
rect 4673 -834 4773 -802
rect 4829 -834 4929 -802
rect 4985 -834 5085 -802
rect 5141 -834 5241 -802
rect 5407 -834 5507 -802
rect 5563 -834 5663 -802
<< polycont >>
rect 135 1783 169 1817
rect 230 1783 264 1817
rect 325 1783 359 1817
rect 557 1783 591 1817
rect 651 1783 685 1817
rect 773 1783 807 1817
rect 867 1783 901 1817
rect 989 1783 1023 1817
rect 1084 1783 1118 1817
rect 1179 1783 1213 1817
rect 1487 1783 1521 1817
rect 1555 1783 1589 1817
rect 1677 1783 1711 1817
rect 1772 1783 1806 1817
rect 1867 1783 1901 1817
rect 1989 1783 2023 1817
rect 2084 1783 2118 1817
rect 2179 1783 2213 1817
rect 2301 1783 2335 1817
rect 2369 1783 2403 1817
rect 2533 1783 2567 1817
rect 2601 1783 2635 1817
rect 2799 1783 2833 1817
rect 2867 1783 2901 1817
rect 2989 1783 3023 1817
rect 3057 1783 3091 1817
rect 105 246 139 280
rect 174 246 208 280
rect 243 246 277 280
rect 312 246 346 280
rect 381 246 415 280
rect 450 246 484 280
rect 519 246 553 280
rect 587 246 621 280
rect 655 246 689 280
rect 723 246 757 280
rect 791 246 825 280
rect 859 246 893 280
rect 927 246 961 280
rect 995 246 1029 280
rect 1063 246 1097 280
rect 1185 246 1219 280
rect 1279 246 1313 280
rect 1401 246 1435 280
rect 1470 246 1504 280
rect 1539 246 1573 280
rect 1608 246 1642 280
rect 1677 246 1711 280
rect 1746 246 1780 280
rect 1815 246 1849 280
rect 1883 246 1917 280
rect 1951 246 1985 280
rect 2019 246 2053 280
rect 2087 246 2121 280
rect 2155 246 2189 280
rect 2223 246 2257 280
rect 2291 246 2325 280
rect 2359 246 2393 280
rect 2481 246 2515 280
rect 2556 246 2590 280
rect 2631 246 2665 280
rect 2705 246 2739 280
rect 2779 246 2813 280
rect 2853 246 2887 280
rect 2927 246 2961 280
rect 3001 246 3035 280
rect 3075 246 3109 280
rect 3149 246 3183 280
rect 3223 246 3257 280
rect 3455 246 3489 280
rect 3549 246 3583 280
rect 3781 246 3815 280
rect 3875 246 3909 280
rect 4107 246 4141 280
rect 4201 246 4235 280
rect 4433 258 4467 292
rect 4508 258 4542 292
rect 4583 258 4617 292
rect 4657 258 4691 292
rect 4731 258 4765 292
rect 4805 258 4839 292
rect 4879 258 4913 292
rect 4953 258 4987 292
rect 5027 258 5061 292
rect 5101 258 5135 292
rect 5175 258 5209 292
rect 5389 246 5423 280
rect 5457 246 5491 280
rect 5579 246 5613 280
rect 5647 246 5681 280
rect 4433 -154 4467 -120
rect 4567 -154 4601 -120
rect 4689 -154 4723 -120
rect 4784 -154 4818 -120
rect 4879 -154 4913 -120
rect 5001 -154 5035 -120
rect 5096 -154 5130 -120
rect 5191 -154 5225 -120
<< locali >>
rect 67 2947 80 2981
rect 135 2947 153 2981
rect 203 2947 226 2981
rect 271 2947 299 2981
rect 339 2947 372 2981
rect 407 2947 441 2981
rect 479 2947 509 2981
rect 552 2947 577 2981
rect 625 2947 645 2981
rect 698 2947 713 2981
rect 771 2947 781 2981
rect 844 2947 849 2981
rect 951 2947 956 2981
rect 1019 2947 1029 2981
rect 1087 2947 1102 2981
rect 1155 2947 1175 2981
rect 1223 2947 1248 2981
rect 1291 2947 1321 2981
rect 1359 2947 1393 2981
rect 1428 2947 1461 2981
rect 1501 2947 1529 2981
rect 1574 2947 1597 2981
rect 1647 2947 1665 2981
rect 1720 2947 1733 2981
rect 1793 2947 1801 2981
rect 1866 2947 1869 2981
rect 1903 2947 1905 2981
rect 1971 2947 1978 2981
rect 2039 2947 2051 2981
rect 2107 2947 2124 2981
rect 2175 2947 2197 2981
rect 2243 2947 2270 2981
rect 2311 2947 2343 2981
rect 2379 2947 2413 2981
rect 2450 2947 2481 2981
rect 2523 2947 2549 2981
rect 2596 2947 2617 2981
rect 2669 2947 2685 2981
rect 2742 2947 2753 2981
rect 2815 2947 2821 2981
rect 2888 2947 2889 2981
rect 2923 2947 2927 2981
rect 2991 2947 3000 2981
rect 3059 2947 3072 2981
rect 3127 2947 3144 2981
rect 3195 2947 3216 2981
rect 3263 2947 3288 2981
rect 3331 2947 3360 2981
rect 3399 2947 3432 2981
rect 3467 2947 3501 2981
rect 3538 2947 3569 2981
rect 3610 2947 3637 2981
rect 3682 2947 3705 2981
rect 3754 2947 3773 2981
rect 3826 2947 3841 2981
rect 3898 2947 3936 2981
rect 3970 2947 3976 2981
rect 74 2795 108 2819
rect 74 2727 108 2742
rect 74 2659 108 2665
rect 74 2622 108 2625
rect 74 2544 108 2557
rect 74 2466 108 2489
rect 74 2388 108 2421
rect 74 2319 108 2353
rect 74 2251 108 2276
rect 74 2183 108 2198
rect 74 2115 108 2120
rect 74 2076 108 2081
rect 74 1998 108 2013
rect 74 1920 108 1945
rect 74 1861 108 1877
rect 230 2795 264 2811
rect 230 2736 264 2761
rect 230 2661 264 2693
rect 230 2591 264 2625
rect 230 2523 264 2552
rect 230 2455 264 2477
rect 230 2387 264 2402
rect 230 2319 264 2327
rect 230 2251 264 2252
rect 230 2211 264 2217
rect 230 2135 264 2149
rect 230 2059 264 2081
rect 230 1983 264 2013
rect 230 1911 264 1945
rect 230 1861 264 1873
rect 386 2795 420 2819
rect 386 2727 420 2745
rect 386 2659 420 2671
rect 386 2591 420 2597
rect 386 2483 420 2489
rect 386 2409 420 2421
rect 386 2335 420 2353
rect 386 2261 420 2285
rect 386 2187 420 2217
rect 386 2115 420 2149
rect 386 2047 420 2079
rect 386 1979 420 2005
rect 386 1911 420 1945
rect 386 1861 420 1877
rect 496 2795 530 2811
rect 496 2736 530 2761
rect 496 2661 530 2693
rect 496 2591 530 2625
rect 496 2523 530 2552
rect 496 2455 530 2477
rect 496 2387 530 2402
rect 496 2319 530 2327
rect 496 2251 530 2252
rect 496 2211 530 2217
rect 496 2135 530 2149
rect 496 2059 530 2081
rect 496 1983 530 2013
rect 496 1911 530 1945
rect 496 1861 530 1873
rect 712 2795 746 2811
rect 712 2736 746 2761
rect 712 2661 746 2693
rect 712 2591 746 2625
rect 712 2523 746 2552
rect 712 2455 746 2477
rect 712 2387 746 2402
rect 712 2319 746 2327
rect 712 2251 746 2252
rect 712 2211 746 2217
rect 712 2135 746 2149
rect 712 2059 746 2081
rect 712 1983 746 2013
rect 712 1911 746 1945
rect 712 1861 746 1873
rect 928 2795 962 2811
rect 928 2736 962 2761
rect 928 2661 962 2693
rect 928 2591 962 2625
rect 928 2523 962 2552
rect 928 2455 962 2477
rect 928 2387 962 2402
rect 928 2319 962 2327
rect 928 2251 962 2252
rect 928 2211 962 2217
rect 928 2135 962 2149
rect 928 2059 962 2081
rect 928 1983 962 2013
rect 928 1911 962 1945
rect 928 1861 962 1873
rect 1084 2795 1118 2819
rect 1084 2727 1118 2745
rect 1084 2659 1118 2671
rect 1084 2591 1118 2597
rect 1084 2483 1118 2489
rect 1084 2409 1118 2421
rect 1084 2335 1118 2353
rect 1084 2261 1118 2285
rect 1084 2187 1118 2217
rect 1084 2115 1118 2149
rect 1084 2047 1118 2078
rect 1084 1979 1118 2003
rect 1084 1911 1118 1945
rect 1084 1861 1118 1877
rect 1240 2795 1274 2811
rect 1240 2736 1274 2761
rect 1240 2661 1274 2693
rect 1240 2591 1274 2625
rect 1240 2523 1274 2552
rect 1240 2455 1274 2477
rect 1240 2387 1274 2402
rect 1240 2319 1274 2327
rect 1240 2251 1274 2252
rect 1240 2211 1274 2217
rect 1240 2135 1274 2149
rect 1240 2059 1274 2081
rect 1240 1983 1274 2013
rect 1240 1911 1274 1945
rect 1240 1861 1274 1873
rect 1400 2795 1434 2819
rect 1400 2727 1434 2747
rect 1400 2659 1434 2675
rect 1400 2591 1434 2603
rect 1400 2523 1434 2530
rect 1400 2455 1434 2457
rect 1400 2418 1434 2421
rect 1400 2345 1434 2353
rect 1400 2272 1434 2285
rect 1400 2199 1434 2217
rect 1400 2126 1434 2149
rect 1400 2053 1434 2081
rect 1400 1980 1434 2013
rect 1400 1911 1434 1945
rect 1400 1861 1434 1873
rect 1616 2795 1650 2819
rect 1616 2727 1650 2747
rect 1616 2659 1650 2675
rect 1616 2591 1650 2603
rect 1616 2523 1650 2530
rect 1616 2455 1650 2457
rect 1616 2418 1650 2421
rect 1616 2345 1650 2353
rect 1616 2272 1650 2285
rect 1616 2199 1650 2217
rect 1616 2126 1650 2149
rect 1616 2053 1650 2081
rect 1616 1980 1650 2013
rect 1616 1911 1650 1945
rect 1616 1861 1650 1873
rect 1772 2795 1806 2811
rect 1772 2736 1806 2761
rect 1772 2661 1806 2693
rect 1772 2591 1806 2625
rect 1772 2523 1806 2552
rect 1772 2455 1806 2477
rect 1772 2387 1806 2402
rect 1772 2319 1806 2327
rect 1772 2251 1806 2252
rect 1772 2211 1806 2217
rect 1772 2135 1806 2149
rect 1772 2059 1806 2081
rect 1772 1983 1806 2013
rect 1772 1911 1806 1945
rect 1772 1861 1806 1873
rect 1928 2795 1962 2819
rect 1928 2727 1962 2747
rect 1928 2659 1962 2675
rect 1928 2591 1962 2603
rect 1928 2523 1962 2530
rect 1928 2455 1962 2457
rect 1928 2418 1962 2421
rect 1928 2345 1962 2353
rect 1928 2272 1962 2285
rect 1928 2199 1962 2217
rect 1928 2126 1962 2149
rect 1928 2053 1962 2081
rect 1928 1980 1962 2013
rect 1928 1911 1962 1945
rect 1928 1861 1962 1873
rect 2084 2795 2118 2811
rect 2084 2736 2118 2761
rect 2084 2661 2118 2693
rect 2084 2591 2118 2625
rect 2084 2523 2118 2552
rect 2084 2455 2118 2477
rect 2084 2387 2118 2402
rect 2084 2319 2118 2327
rect 2084 2251 2118 2252
rect 2084 2211 2118 2217
rect 2084 2135 2118 2149
rect 2084 2059 2118 2081
rect 2084 1983 2118 2013
rect 2084 1911 2118 1945
rect 2084 1861 2118 1873
rect 2240 2795 2274 2819
rect 2240 2727 2274 2747
rect 2240 2659 2274 2675
rect 2240 2591 2274 2603
rect 2240 2523 2274 2530
rect 2240 2455 2274 2457
rect 2240 2418 2274 2421
rect 2240 2345 2274 2353
rect 2240 2272 2274 2285
rect 2240 2199 2274 2217
rect 2240 2126 2274 2149
rect 2240 2053 2274 2081
rect 2240 1980 2274 2013
rect 2240 1911 2274 1945
rect 2240 1861 2274 1873
rect 2396 2795 2430 2811
rect 2396 2736 2430 2761
rect 2396 2661 2430 2693
rect 2396 2591 2430 2625
rect 2396 2523 2430 2552
rect 2396 2455 2430 2477
rect 2772 2795 2806 2811
rect 2772 2736 2806 2761
rect 2772 2659 2806 2693
rect 2772 2591 2806 2624
rect 2772 2523 2806 2546
rect 2772 2455 2806 2468
rect 2396 2387 2430 2402
rect 2396 2319 2430 2327
rect 2396 2251 2430 2252
rect 2396 2211 2430 2217
rect 2396 2135 2430 2149
rect 2396 2059 2430 2081
rect 2396 1983 2430 2013
rect 2396 1911 2430 1945
rect 2396 1861 2430 1873
rect 2506 2387 2540 2403
rect 2506 2319 2540 2332
rect 2506 2281 2540 2285
rect 2506 2196 2540 2217
rect 2506 2115 2540 2149
rect 2506 2047 2540 2077
rect 2506 1979 2540 1992
rect 2506 1941 2540 1945
rect 2506 1861 2540 1877
rect 2662 2387 2696 2403
rect 2662 2319 2696 2332
rect 2662 2281 2696 2285
rect 2662 2196 2696 2217
rect 2662 2115 2696 2149
rect 2662 2047 2696 2077
rect 2662 1979 2696 1992
rect 2662 1941 2696 1945
rect 2662 1861 2696 1877
rect 2772 2387 2806 2390
rect 2772 2346 2806 2353
rect 2772 2267 2806 2285
rect 2772 2188 2806 2217
rect 2772 2115 2806 2149
rect 2772 2047 2806 2075
rect 2772 1979 2806 1996
rect 2772 1911 2806 1945
rect 2772 1861 2806 1877
rect 2928 2795 2962 2819
rect 2928 2727 2962 2742
rect 2928 2659 2962 2665
rect 2928 2621 2962 2625
rect 2928 2543 2962 2557
rect 2928 2465 2962 2489
rect 2928 2387 2962 2421
rect 2928 2319 2962 2353
rect 2928 2251 2962 2275
rect 2928 2183 2962 2197
rect 2928 2115 2962 2119
rect 2928 2075 2962 2081
rect 2928 1997 2962 2013
rect 2928 1911 2962 1945
rect 2928 1861 2962 1877
rect 3084 2795 3118 2811
rect 3084 2736 3118 2761
rect 3084 2661 3118 2693
rect 3084 2591 3118 2625
rect 3084 2523 3118 2552
rect 3084 2455 3118 2477
rect 3492 2405 3530 2439
rect 3084 2387 3118 2402
rect 3084 2319 3118 2327
rect 3430 2262 3468 2296
rect 3646 2287 3680 2325
rect 3791 2299 3825 2337
rect 3894 2286 3928 2324
rect 3084 2251 3118 2252
rect 3084 2211 3118 2217
rect 3084 2136 3118 2149
rect 3084 2060 3118 2081
rect 3084 1984 3118 2013
rect 3084 1911 3118 1945
rect 3084 1861 3118 1877
rect 119 1783 135 1817
rect 171 1783 230 1817
rect 265 1783 324 1817
rect 359 1783 375 1817
rect 541 1783 557 1817
rect 612 1783 650 1817
rect 685 1783 701 1817
rect 757 1783 773 1817
rect 818 1783 856 1817
rect 901 1783 917 1817
rect 973 1783 985 1817
rect 1023 1783 1084 1817
rect 1118 1783 1179 1817
rect 1217 1783 1229 1817
rect 1441 1783 1479 1817
rect 1521 1783 1555 1817
rect 1589 1783 1605 1817
rect 1661 1783 1673 1817
rect 1711 1783 1767 1817
rect 1806 1783 1860 1817
rect 1901 1783 1917 1817
rect 1973 1783 1989 1817
rect 2026 1783 2084 1817
rect 2120 1783 2179 1817
rect 2213 1783 2229 1817
rect 2285 1783 2301 1817
rect 2340 1783 2369 1817
rect 2412 1783 2419 1817
rect 2567 1783 2582 1817
rect 2635 1783 2651 1817
rect 2783 1783 2795 1817
rect 2833 1783 2867 1817
rect 2901 1783 2917 1817
rect 2973 1783 2987 1817
rect 3023 1783 3057 1817
rect 3093 1783 3107 1817
rect 89 246 105 280
rect 146 246 174 280
rect 223 246 243 280
rect 300 246 312 280
rect 377 246 381 280
rect 415 246 420 280
rect 484 246 497 280
rect 553 246 574 280
rect 621 246 651 280
rect 689 246 723 280
rect 762 246 791 280
rect 839 246 859 280
rect 916 246 927 280
rect 992 246 995 280
rect 1029 246 1034 280
rect 1097 246 1113 280
rect 1169 246 1185 280
rect 1232 246 1270 280
rect 1313 246 1329 280
rect 1385 246 1401 280
rect 1449 246 1470 280
rect 1526 246 1539 280
rect 1603 246 1608 280
rect 1642 246 1646 280
rect 1711 246 1723 280
rect 1780 246 1800 280
rect 1849 246 1877 280
rect 1917 246 1951 280
rect 1988 246 2019 280
rect 2065 246 2087 280
rect 2142 246 2155 280
rect 2219 246 2223 280
rect 2257 246 2261 280
rect 2325 246 2337 280
rect 2393 246 2409 280
rect 2465 246 2481 280
rect 2541 246 2556 280
rect 2619 246 2631 280
rect 2697 246 2705 280
rect 2739 246 2741 280
rect 2775 246 2779 280
rect 2813 246 2819 280
rect 2887 246 2896 280
rect 2961 246 2973 280
rect 3035 246 3050 280
rect 3109 246 3127 280
rect 3183 246 3204 280
rect 3257 246 3273 280
rect 3439 246 3455 280
rect 3507 246 3545 280
rect 3583 246 3599 280
rect 3765 246 3781 280
rect 3833 246 3871 280
rect 3909 246 3925 280
rect 4091 246 4107 280
rect 4159 246 4197 280
rect 4235 246 4251 280
rect 4417 258 4433 292
rect 4467 285 4508 292
rect 4542 285 4583 292
rect 4617 285 4657 292
rect 4691 285 4731 292
rect 4765 285 4805 292
rect 4839 285 4879 292
rect 4913 285 4953 292
rect 4987 285 5027 292
rect 5061 285 5101 292
rect 5135 285 5175 292
rect 4467 258 4489 285
rect 4542 258 4562 285
rect 4617 258 4635 285
rect 4691 258 4708 285
rect 4765 258 4781 285
rect 4839 258 4854 285
rect 4913 258 4926 285
rect 4987 258 4998 285
rect 5061 258 5070 285
rect 5135 258 5142 285
rect 5209 258 5225 292
rect 4523 251 4562 258
rect 4596 251 4635 258
rect 4669 251 4708 258
rect 4742 251 4781 258
rect 4815 251 4854 258
rect 4888 251 4926 258
rect 4960 251 4998 258
rect 5032 251 5070 258
rect 5104 251 5142 258
rect 5423 246 5433 280
rect 5491 246 5507 280
rect 5563 246 5577 280
rect 5613 246 5647 280
rect 5683 246 5697 280
rect 4372 201 4406 217
rect 44 128 78 162
rect 44 60 78 88
rect 44 -8 78 14
rect 44 -76 78 -60
rect 44 -144 78 -134
rect 44 -212 78 -208
rect 44 -248 78 -246
rect 44 -322 78 -314
rect 44 -395 78 -382
rect 44 -468 78 -450
rect 44 -541 78 -518
rect 44 -614 78 -586
rect 44 -687 78 -654
rect 44 -756 78 -722
rect 44 -806 78 -794
rect 260 128 294 162
rect 260 60 294 87
rect 260 -8 294 12
rect 260 -76 294 -63
rect 260 -144 294 -138
rect 260 -179 294 -178
rect 260 -254 294 -246
rect 260 -329 294 -314
rect 260 -404 294 -382
rect 260 -479 294 -450
rect 260 -552 294 -518
rect 260 -620 294 -588
rect 260 -688 294 -662
rect 260 -756 294 -722
rect 260 -806 294 -790
rect 476 128 510 144
rect 476 64 510 94
rect 476 -8 510 26
rect 476 -76 510 -45
rect 476 -144 510 -120
rect 476 -212 510 -195
rect 476 -280 510 -270
rect 476 -348 510 -345
rect 476 -386 510 -382
rect 476 -461 510 -450
rect 476 -536 510 -518
rect 476 -611 510 -586
rect 476 -686 510 -654
rect 476 -756 510 -722
rect 476 -806 510 -794
rect 692 128 726 162
rect 692 60 726 87
rect 692 -8 726 12
rect 692 -76 726 -63
rect 692 -144 726 -138
rect 692 -179 726 -178
rect 692 -254 726 -246
rect 692 -329 726 -314
rect 692 -404 726 -382
rect 692 -479 726 -450
rect 692 -552 726 -518
rect 692 -620 726 -588
rect 692 -688 726 -662
rect 692 -756 726 -722
rect 692 -806 726 -790
rect 908 128 942 144
rect 908 64 942 94
rect 908 -8 942 26
rect 908 -76 942 -45
rect 908 -144 942 -120
rect 908 -212 942 -195
rect 908 -280 942 -270
rect 908 -348 942 -345
rect 908 -386 942 -382
rect 908 -461 942 -450
rect 908 -536 942 -518
rect 908 -611 942 -586
rect 908 -686 942 -654
rect 908 -756 942 -722
rect 908 -806 942 -794
rect 1124 128 1158 162
rect 1124 60 1158 87
rect 1124 -8 1158 12
rect 1124 -76 1158 -63
rect 1124 -144 1158 -138
rect 1124 -179 1158 -178
rect 1124 -254 1158 -246
rect 1124 -329 1158 -314
rect 1124 -404 1158 -382
rect 1124 -479 1158 -450
rect 1124 -552 1158 -518
rect 1124 -620 1158 -588
rect 1124 -688 1158 -662
rect 1124 -756 1158 -722
rect 1124 -806 1158 -790
rect 1340 128 1374 144
rect 1340 64 1374 94
rect 1340 -8 1374 26
rect 1340 -76 1374 -45
rect 1340 -144 1374 -120
rect 1340 -212 1374 -195
rect 1340 -280 1374 -270
rect 1340 -348 1374 -345
rect 1340 -386 1374 -382
rect 1340 -461 1374 -450
rect 1340 -536 1374 -518
rect 1340 -611 1374 -586
rect 1340 -686 1374 -654
rect 1340 -756 1374 -722
rect 1340 -806 1374 -794
rect 1556 128 1590 162
rect 1556 60 1590 87
rect 1556 -8 1590 12
rect 1556 -76 1590 -63
rect 1556 -144 1590 -138
rect 1556 -179 1590 -178
rect 1556 -254 1590 -246
rect 1556 -329 1590 -314
rect 1556 -404 1590 -382
rect 1556 -479 1590 -450
rect 1556 -552 1590 -518
rect 1556 -620 1590 -588
rect 1556 -688 1590 -662
rect 1556 -756 1590 -722
rect 1556 -806 1590 -790
rect 1772 128 1806 144
rect 1772 64 1806 94
rect 1772 -8 1806 26
rect 1772 -76 1806 -45
rect 1772 -144 1806 -120
rect 1772 -212 1806 -195
rect 1772 -280 1806 -270
rect 1772 -348 1806 -345
rect 1772 -386 1806 -382
rect 1772 -461 1806 -450
rect 1772 -536 1806 -518
rect 1772 -611 1806 -586
rect 1772 -686 1806 -654
rect 1772 -756 1806 -722
rect 1772 -806 1806 -794
rect 1988 128 2022 162
rect 1988 60 2022 87
rect 1988 -8 2022 12
rect 1988 -76 2022 -63
rect 1988 -144 2022 -138
rect 1988 -179 2022 -178
rect 1988 -254 2022 -246
rect 1988 -329 2022 -314
rect 1988 -404 2022 -382
rect 1988 -479 2022 -450
rect 1988 -552 2022 -518
rect 1988 -620 2022 -588
rect 1988 -688 2022 -662
rect 1988 -756 2022 -722
rect 1988 -806 2022 -790
rect 2204 128 2238 144
rect 2204 64 2238 94
rect 2204 -8 2238 26
rect 2204 -76 2238 -45
rect 2204 -144 2238 -120
rect 2204 -212 2238 -195
rect 2204 -280 2238 -270
rect 2204 -348 2238 -345
rect 2204 -386 2238 -382
rect 2204 -461 2238 -450
rect 2204 -536 2238 -518
rect 2204 -611 2238 -586
rect 2204 -686 2238 -654
rect 2204 -756 2238 -722
rect 2204 -806 2238 -794
rect 2420 128 2454 162
rect 2420 60 2454 87
rect 2420 -8 2454 12
rect 2420 -76 2454 -63
rect 2420 -144 2454 -138
rect 2420 -179 2454 -178
rect 2420 -254 2454 -246
rect 2420 -329 2454 -314
rect 2420 -404 2454 -382
rect 2420 -479 2454 -450
rect 2420 -552 2454 -518
rect 2420 -620 2454 -588
rect 2420 -688 2454 -662
rect 2420 -756 2454 -722
rect 2420 -806 2454 -790
rect 2636 128 2670 144
rect 2636 64 2670 94
rect 2636 -8 2670 26
rect 2636 -76 2670 -45
rect 2636 -144 2670 -120
rect 2636 -212 2670 -195
rect 2636 -280 2670 -270
rect 2636 -348 2670 -345
rect 2636 -386 2670 -382
rect 2636 -461 2670 -450
rect 2636 -536 2670 -518
rect 2636 -611 2670 -586
rect 2636 -686 2670 -654
rect 2636 -756 2670 -722
rect 2636 -806 2670 -794
rect 2852 128 2886 162
rect 2852 60 2886 87
rect 2852 -8 2886 12
rect 2852 -76 2886 -63
rect 2852 -144 2886 -138
rect 2852 -179 2886 -178
rect 2852 -254 2886 -246
rect 2852 -329 2886 -314
rect 2852 -404 2886 -382
rect 2852 -479 2886 -450
rect 2852 -552 2886 -518
rect 2852 -620 2886 -588
rect 2852 -688 2886 -662
rect 2852 -756 2886 -722
rect 2852 -806 2886 -790
rect 3068 128 3102 144
rect 3068 64 3102 94
rect 3068 -8 3102 26
rect 3068 -76 3102 -45
rect 3068 -144 3102 -120
rect 3068 -212 3102 -195
rect 3068 -280 3102 -270
rect 3068 -348 3102 -345
rect 3068 -386 3102 -382
rect 3068 -461 3102 -450
rect 3068 -536 3102 -518
rect 3068 -611 3102 -586
rect 3068 -686 3102 -654
rect 3068 -756 3102 -722
rect 3068 -806 3102 -794
rect 3284 128 3318 162
rect 3284 60 3318 87
rect 3284 -8 3318 12
rect 3284 -76 3318 -63
rect 3284 -144 3318 -138
rect 3284 -179 3318 -178
rect 3284 -254 3318 -246
rect 3284 -329 3318 -314
rect 3284 -404 3318 -382
rect 3284 -479 3318 -450
rect 3284 -552 3318 -518
rect 3284 -620 3318 -588
rect 3284 -688 3318 -662
rect 3284 -756 3318 -722
rect 3284 -806 3318 -790
rect 3394 128 3428 162
rect 3394 60 3428 87
rect 3394 -8 3428 12
rect 3394 -76 3428 -63
rect 3394 -144 3428 -138
rect 3394 -179 3428 -178
rect 3394 -254 3428 -246
rect 3394 -329 3428 -314
rect 3394 -404 3428 -382
rect 3394 -479 3428 -450
rect 3394 -552 3428 -518
rect 3394 -620 3428 -588
rect 3394 -688 3428 -662
rect 3394 -756 3428 -722
rect 3394 -806 3428 -790
rect 3610 128 3644 144
rect 3610 64 3644 94
rect 3610 -8 3644 26
rect 3610 -76 3644 -45
rect 3610 -144 3644 -120
rect 3610 -212 3644 -195
rect 3610 -280 3644 -270
rect 3610 -348 3644 -345
rect 3610 -386 3644 -382
rect 3610 -461 3644 -450
rect 3610 -536 3644 -518
rect 3610 -611 3644 -586
rect 3610 -686 3644 -654
rect 3610 -756 3644 -722
rect 3610 -806 3644 -794
rect 3720 128 3754 144
rect 3720 64 3754 94
rect 3720 -8 3754 26
rect 3720 -76 3754 -45
rect 3720 -144 3754 -120
rect 3720 -212 3754 -195
rect 3720 -280 3754 -270
rect 3720 -348 3754 -345
rect 3720 -386 3754 -382
rect 3720 -461 3754 -450
rect 3720 -536 3754 -518
rect 3720 -611 3754 -586
rect 3720 -686 3754 -654
rect 3720 -756 3754 -722
rect 3720 -806 3754 -794
rect 3936 128 3970 144
rect 3936 64 3970 94
rect 3936 -8 3970 26
rect 3936 -76 3970 -45
rect 3936 -144 3970 -120
rect 3936 -212 3970 -195
rect 3936 -280 3970 -270
rect 3936 -348 3970 -345
rect 3936 -386 3970 -382
rect 3936 -461 3970 -450
rect 3936 -536 3970 -518
rect 3936 -611 3970 -586
rect 3936 -686 3970 -654
rect 3936 -756 3970 -722
rect 3936 -806 3970 -794
rect 4046 128 4080 144
rect 4046 64 4080 94
rect 4046 -8 4080 26
rect 4046 -76 4080 -45
rect 4046 -144 4080 -120
rect 4046 -212 4080 -195
rect 4046 -280 4080 -270
rect 4046 -348 4080 -345
rect 4046 -386 4080 -382
rect 4046 -461 4080 -450
rect 4046 -536 4080 -518
rect 4046 -611 4080 -586
rect 4046 -686 4080 -654
rect 4046 -756 4080 -722
rect 4046 -806 4080 -794
rect 4262 128 4296 144
rect 4262 64 4296 94
rect 4262 -8 4296 26
rect 4372 133 4406 162
rect 4372 65 4406 90
rect 4588 201 4622 217
rect 4588 133 4622 167
rect 4588 65 4622 99
rect 4372 15 4406 31
rect 4586 31 4588 41
rect 4804 201 4838 217
rect 4804 133 4838 162
rect 4804 65 4838 90
rect 4622 31 4624 41
rect 4586 7 4624 31
rect 5020 201 5054 217
rect 5020 133 5054 167
rect 5020 65 5054 99
rect 4804 15 4838 31
rect 5018 31 5020 41
rect 5236 201 5270 217
rect 5236 133 5270 162
rect 5236 65 5270 90
rect 5054 31 5056 41
rect 5018 7 5056 31
rect 5236 15 5270 31
rect 5362 128 5396 144
rect 5362 60 5396 94
rect 5362 19 5396 26
rect 4262 -76 4296 -45
rect 5362 -56 5396 -42
rect 4719 -120 4777 -119
rect 4811 -120 4868 -119
rect 4262 -144 4296 -120
rect 4417 -154 4433 -120
rect 4467 -154 4471 -120
rect 4505 -154 4543 -120
rect 4601 -154 4617 -120
rect 4673 -153 4685 -120
rect 4723 -153 4777 -120
rect 4818 -153 4868 -120
rect 4673 -154 4689 -153
rect 4723 -154 4784 -153
rect 4818 -154 4879 -153
rect 4913 -154 4929 -120
rect 4985 -154 4997 -120
rect 5035 -154 5081 -120
rect 5130 -154 5165 -120
rect 5225 -154 5241 -120
rect 5362 -131 5396 -110
rect 4262 -212 4296 -195
rect 5362 -206 5396 -178
rect 4262 -280 4296 -270
rect 4262 -348 4296 -345
rect 4262 -386 4296 -382
rect 4262 -461 4296 -450
rect 4262 -536 4296 -518
rect 4262 -611 4296 -586
rect 4262 -686 4296 -654
rect 4262 -756 4296 -722
rect 4262 -806 4296 -794
rect 4372 -339 4406 -314
rect 4372 -415 4406 -382
rect 4372 -484 4406 -450
rect 4372 -552 4406 -525
rect 4372 -620 4406 -601
rect 4372 -688 4406 -677
rect 4372 -756 4406 -722
rect 4372 -806 4406 -790
rect 4628 -280 4662 -264
rect 4628 -348 4662 -314
rect 4628 -416 4662 -415
rect 4628 -456 4662 -450
rect 4628 -532 4662 -518
rect 4628 -608 4662 -586
rect 4628 -684 4662 -654
rect 4628 -756 4662 -722
rect 4628 -806 4662 -794
rect 4784 -276 4818 -264
rect 4784 -348 4818 -314
rect 4784 -416 4818 -385
rect 4784 -484 4818 -461
rect 4784 -552 4818 -537
rect 4784 -620 4818 -613
rect 4784 -655 4818 -654
rect 4784 -756 4818 -722
rect 4784 -806 4818 -790
rect 4940 -280 4974 -264
rect 4940 -348 4974 -314
rect 4940 -416 4974 -415
rect 4940 -456 4974 -450
rect 4940 -532 4974 -518
rect 4940 -608 4974 -586
rect 4940 -684 4974 -654
rect 4940 -756 4974 -722
rect 4940 -806 4974 -794
rect 5096 -276 5130 -264
rect 5096 -348 5130 -314
rect 5096 -416 5130 -385
rect 5096 -484 5130 -461
rect 5096 -552 5130 -537
rect 5096 -620 5130 -613
rect 5096 -655 5130 -654
rect 5096 -756 5130 -722
rect 5096 -806 5130 -790
rect 5252 -280 5286 -264
rect 5252 -348 5286 -314
rect 5252 -416 5286 -415
rect 5252 -456 5286 -450
rect 5252 -532 5286 -518
rect 5252 -608 5286 -586
rect 5252 -684 5286 -654
rect 5252 -756 5286 -722
rect 5252 -806 5286 -794
rect 5362 -280 5396 -246
rect 5362 -348 5396 -315
rect 5362 -416 5396 -390
rect 5362 -484 5396 -465
rect 5362 -552 5396 -540
rect 5362 -620 5396 -616
rect 5362 -688 5396 -654
rect 5362 -756 5396 -722
rect 5362 -806 5396 -790
rect 5518 128 5552 144
rect 5518 60 5552 94
rect 5518 19 5552 26
rect 5518 -58 5552 -42
rect 5518 -136 5552 -110
rect 5518 -212 5552 -178
rect 5518 -280 5552 -248
rect 5518 -348 5552 -326
rect 5518 -416 5552 -404
rect 5518 -484 5552 -482
rect 5518 -526 5552 -518
rect 5518 -604 5552 -586
rect 5518 -682 5552 -654
rect 5518 -756 5552 -722
rect 5518 -806 5552 -794
rect 5674 128 5708 144
rect 5674 75 5675 94
rect 5674 60 5709 75
rect 5708 33 5709 60
rect 5674 -1 5675 26
rect 5674 -8 5709 -1
rect 5708 -42 5709 -8
rect 5674 -43 5709 -42
rect 5674 -76 5675 -43
rect 5708 -110 5709 -77
rect 5674 -120 5709 -110
rect 5674 -144 5675 -120
rect 5708 -178 5709 -154
rect 5674 -197 5709 -178
rect 5674 -212 5675 -197
rect 5708 -246 5709 -231
rect 5674 -274 5709 -246
rect 5674 -280 5675 -274
rect 5708 -314 5709 -308
rect 5674 -348 5709 -314
rect 5708 -351 5709 -348
rect 5674 -385 5675 -382
rect 5674 -416 5709 -385
rect 5708 -428 5709 -416
rect 5674 -462 5675 -450
rect 5674 -484 5709 -462
rect 5708 -505 5709 -484
rect 5674 -539 5675 -518
rect 5674 -552 5709 -539
rect 5708 -582 5709 -552
rect 5674 -616 5675 -586
rect 5674 -620 5708 -616
rect 5674 -688 5708 -654
rect 5674 -756 5708 -722
rect 5674 -806 5708 -790
rect 125 -912 140 -878
rect 194 -912 213 -878
rect 263 -912 286 -878
rect 332 -912 359 -878
rect 401 -912 432 -878
rect 470 -912 505 -878
rect 539 -912 574 -878
rect 612 -912 643 -878
rect 685 -912 712 -878
rect 758 -912 781 -878
rect 831 -912 850 -878
rect 904 -912 919 -878
rect 977 -912 988 -878
rect 1050 -912 1057 -878
rect 1123 -912 1126 -878
rect 1160 -912 1162 -878
rect 1229 -912 1235 -878
rect 1298 -912 1308 -878
rect 1367 -912 1381 -878
rect 1436 -912 1454 -878
rect 1505 -912 1527 -878
rect 1574 -912 1600 -878
rect 1643 -912 1673 -878
rect 1712 -912 1746 -878
rect 1781 -912 1816 -878
rect 1853 -912 1885 -878
rect 1926 -912 1954 -878
rect 1999 -912 2023 -878
rect 2072 -912 2092 -878
rect 2145 -912 2161 -878
rect 2218 -912 2230 -878
rect 2291 -912 2299 -878
rect 2364 -912 2368 -878
rect 2402 -912 2403 -878
rect 2471 -912 2476 -878
rect 2539 -912 2549 -878
rect 2607 -912 2622 -878
rect 2675 -912 2695 -878
rect 2743 -912 2768 -878
rect 2811 -912 2841 -878
rect 2879 -912 2913 -878
rect 2948 -912 2981 -878
rect 3021 -912 3049 -878
rect 3094 -912 3117 -878
rect 3167 -912 3185 -878
rect 3240 -912 3253 -878
rect 3313 -912 3321 -878
rect 3386 -912 3389 -878
rect 3423 -912 3425 -878
rect 3491 -912 3498 -878
rect 3559 -912 3570 -878
rect 3627 -912 3642 -878
rect 3695 -912 3714 -878
rect 3763 -912 3786 -878
rect 3831 -912 3858 -878
rect 3899 -912 3930 -878
rect 3967 -912 4001 -878
rect 4036 -912 4069 -878
rect 4108 -912 4137 -878
rect 4180 -912 4205 -878
rect 4252 -912 4273 -878
rect 4324 -912 4341 -878
rect 4396 -912 4409 -878
rect 4468 -912 4477 -878
rect 4540 -912 4545 -878
rect 4612 -912 4613 -878
rect 4647 -912 4650 -878
rect 4715 -912 4722 -878
rect 4783 -912 4794 -878
rect 4851 -912 4866 -878
rect 4919 -912 4938 -878
rect 4987 -912 5010 -878
rect 5055 -912 5082 -878
rect 5123 -912 5154 -878
rect 5191 -912 5225 -878
rect 5260 -912 5293 -878
rect 5332 -912 5361 -878
rect 5404 -912 5429 -878
rect 5476 -912 5497 -878
rect 5548 -912 5565 -878
rect 5620 -912 5633 -878
<< viali >>
rect 80 2947 101 2981
rect 101 2947 114 2981
rect 153 2947 169 2981
rect 169 2947 187 2981
rect 226 2947 237 2981
rect 237 2947 260 2981
rect 299 2947 305 2981
rect 305 2947 333 2981
rect 372 2947 373 2981
rect 373 2947 406 2981
rect 445 2947 475 2981
rect 475 2947 479 2981
rect 518 2947 543 2981
rect 543 2947 552 2981
rect 591 2947 611 2981
rect 611 2947 625 2981
rect 664 2947 679 2981
rect 679 2947 698 2981
rect 737 2947 747 2981
rect 747 2947 771 2981
rect 810 2947 815 2981
rect 815 2947 844 2981
rect 883 2947 917 2981
rect 956 2947 985 2981
rect 985 2947 990 2981
rect 1029 2947 1053 2981
rect 1053 2947 1063 2981
rect 1102 2947 1121 2981
rect 1121 2947 1136 2981
rect 1175 2947 1189 2981
rect 1189 2947 1209 2981
rect 1248 2947 1257 2981
rect 1257 2947 1282 2981
rect 1321 2947 1325 2981
rect 1325 2947 1355 2981
rect 1394 2947 1427 2981
rect 1427 2947 1428 2981
rect 1467 2947 1495 2981
rect 1495 2947 1501 2981
rect 1540 2947 1563 2981
rect 1563 2947 1574 2981
rect 1613 2947 1631 2981
rect 1631 2947 1647 2981
rect 1686 2947 1699 2981
rect 1699 2947 1720 2981
rect 1759 2947 1767 2981
rect 1767 2947 1793 2981
rect 1832 2947 1835 2981
rect 1835 2947 1866 2981
rect 1905 2947 1937 2981
rect 1937 2947 1939 2981
rect 1978 2947 2005 2981
rect 2005 2947 2012 2981
rect 2051 2947 2073 2981
rect 2073 2947 2085 2981
rect 2124 2947 2141 2981
rect 2141 2947 2158 2981
rect 2197 2947 2209 2981
rect 2209 2947 2231 2981
rect 2270 2947 2277 2981
rect 2277 2947 2304 2981
rect 2343 2947 2345 2981
rect 2345 2947 2377 2981
rect 2416 2947 2447 2981
rect 2447 2947 2450 2981
rect 2489 2947 2515 2981
rect 2515 2947 2523 2981
rect 2562 2947 2583 2981
rect 2583 2947 2596 2981
rect 2635 2947 2651 2981
rect 2651 2947 2669 2981
rect 2708 2947 2719 2981
rect 2719 2947 2742 2981
rect 2781 2947 2787 2981
rect 2787 2947 2815 2981
rect 2854 2947 2855 2981
rect 2855 2947 2888 2981
rect 2927 2947 2957 2981
rect 2957 2947 2961 2981
rect 3000 2947 3025 2981
rect 3025 2947 3034 2981
rect 3072 2947 3093 2981
rect 3093 2947 3106 2981
rect 3144 2947 3161 2981
rect 3161 2947 3178 2981
rect 3216 2947 3229 2981
rect 3229 2947 3250 2981
rect 3288 2947 3297 2981
rect 3297 2947 3322 2981
rect 3360 2947 3365 2981
rect 3365 2947 3394 2981
rect 3432 2947 3433 2981
rect 3433 2947 3466 2981
rect 3504 2947 3535 2981
rect 3535 2947 3538 2981
rect 3576 2947 3603 2981
rect 3603 2947 3610 2981
rect 3648 2947 3671 2981
rect 3671 2947 3682 2981
rect 3720 2947 3739 2981
rect 3739 2947 3754 2981
rect 3792 2947 3807 2981
rect 3807 2947 3826 2981
rect 3864 2947 3875 2981
rect 3875 2947 3898 2981
rect 3936 2947 3970 2981
rect 74 2819 108 2853
rect 386 2819 420 2853
rect 74 2761 108 2776
rect 74 2742 108 2761
rect 74 2693 108 2699
rect 74 2665 108 2693
rect 74 2591 108 2622
rect 74 2588 108 2591
rect 74 2523 108 2544
rect 74 2510 108 2523
rect 74 2455 108 2466
rect 74 2432 108 2455
rect 74 2387 108 2388
rect 74 2354 108 2387
rect 74 2285 108 2310
rect 74 2276 108 2285
rect 74 2217 108 2232
rect 74 2198 108 2217
rect 74 2149 108 2154
rect 74 2120 108 2149
rect 74 2047 108 2076
rect 74 2042 108 2047
rect 74 1979 108 1998
rect 74 1964 108 1979
rect 74 1911 108 1920
rect 74 1886 108 1911
rect 230 2727 264 2736
rect 230 2702 264 2727
rect 230 2659 264 2661
rect 230 2627 264 2659
rect 230 2557 264 2586
rect 230 2552 264 2557
rect 230 2489 264 2511
rect 230 2477 264 2489
rect 230 2421 264 2436
rect 230 2402 264 2421
rect 230 2353 264 2361
rect 230 2327 264 2353
rect 230 2285 264 2286
rect 230 2252 264 2285
rect 230 2183 264 2211
rect 230 2177 264 2183
rect 230 2115 264 2135
rect 230 2101 264 2115
rect 230 2047 264 2059
rect 230 2025 264 2047
rect 230 1979 264 1983
rect 230 1949 264 1979
rect 230 1877 264 1907
rect 230 1873 264 1877
rect 1084 2819 1118 2853
rect 386 2761 420 2779
rect 386 2745 420 2761
rect 386 2693 420 2705
rect 386 2671 420 2693
rect 386 2625 420 2631
rect 386 2597 420 2625
rect 386 2523 420 2557
rect 386 2455 420 2483
rect 386 2449 420 2455
rect 386 2387 420 2409
rect 386 2375 420 2387
rect 386 2319 420 2335
rect 386 2301 420 2319
rect 386 2251 420 2261
rect 386 2227 420 2251
rect 386 2183 420 2187
rect 386 2153 420 2183
rect 386 2081 420 2113
rect 386 2079 420 2081
rect 386 2013 420 2039
rect 386 2005 420 2013
rect 496 2727 530 2736
rect 496 2702 530 2727
rect 496 2659 530 2661
rect 496 2627 530 2659
rect 496 2557 530 2586
rect 496 2552 530 2557
rect 496 2489 530 2511
rect 496 2477 530 2489
rect 496 2421 530 2436
rect 496 2402 530 2421
rect 496 2353 530 2361
rect 496 2327 530 2353
rect 496 2285 530 2286
rect 496 2252 530 2285
rect 496 2183 530 2211
rect 496 2177 530 2183
rect 496 2115 530 2135
rect 496 2101 530 2115
rect 496 2047 530 2059
rect 496 2025 530 2047
rect 496 1979 530 1983
rect 496 1949 530 1979
rect 496 1877 530 1907
rect 496 1873 530 1877
rect 712 2727 746 2736
rect 712 2702 746 2727
rect 712 2659 746 2661
rect 712 2627 746 2659
rect 712 2557 746 2586
rect 712 2552 746 2557
rect 712 2489 746 2511
rect 712 2477 746 2489
rect 712 2421 746 2436
rect 712 2402 746 2421
rect 712 2353 746 2361
rect 712 2327 746 2353
rect 712 2285 746 2286
rect 712 2252 746 2285
rect 712 2183 746 2211
rect 712 2177 746 2183
rect 712 2115 746 2135
rect 712 2101 746 2115
rect 712 2047 746 2059
rect 712 2025 746 2047
rect 712 1979 746 1983
rect 712 1949 746 1979
rect 712 1877 746 1907
rect 712 1873 746 1877
rect 928 2727 962 2736
rect 928 2702 962 2727
rect 928 2659 962 2661
rect 928 2627 962 2659
rect 928 2557 962 2586
rect 928 2552 962 2557
rect 928 2489 962 2511
rect 928 2477 962 2489
rect 928 2421 962 2436
rect 928 2402 962 2421
rect 928 2353 962 2361
rect 928 2327 962 2353
rect 928 2285 962 2286
rect 928 2252 962 2285
rect 928 2183 962 2211
rect 928 2177 962 2183
rect 928 2115 962 2135
rect 928 2101 962 2115
rect 928 2047 962 2059
rect 928 2025 962 2047
rect 928 1979 962 1983
rect 928 1949 962 1979
rect 928 1877 962 1907
rect 928 1873 962 1877
rect 1400 2819 1434 2853
rect 1084 2761 1118 2779
rect 1084 2745 1118 2761
rect 1084 2693 1118 2705
rect 1084 2671 1118 2693
rect 1084 2625 1118 2631
rect 1084 2597 1118 2625
rect 1084 2523 1118 2557
rect 1084 2455 1118 2483
rect 1084 2449 1118 2455
rect 1084 2387 1118 2409
rect 1084 2375 1118 2387
rect 1084 2319 1118 2335
rect 1084 2301 1118 2319
rect 1084 2251 1118 2261
rect 1084 2227 1118 2251
rect 1084 2183 1118 2187
rect 1084 2153 1118 2183
rect 1084 2081 1118 2112
rect 1084 2078 1118 2081
rect 1084 2013 1118 2037
rect 1084 2003 1118 2013
rect 1240 2727 1274 2736
rect 1240 2702 1274 2727
rect 1240 2659 1274 2661
rect 1240 2627 1274 2659
rect 1240 2557 1274 2586
rect 1240 2552 1274 2557
rect 1240 2489 1274 2511
rect 1240 2477 1274 2489
rect 1240 2421 1274 2436
rect 1240 2402 1274 2421
rect 1240 2353 1274 2361
rect 1240 2327 1274 2353
rect 1240 2285 1274 2286
rect 1240 2252 1274 2285
rect 1240 2183 1274 2211
rect 1240 2177 1274 2183
rect 1240 2115 1274 2135
rect 1240 2101 1274 2115
rect 1240 2047 1274 2059
rect 1240 2025 1274 2047
rect 1240 1979 1274 1983
rect 1240 1949 1274 1979
rect 1240 1877 1274 1907
rect 1240 1873 1274 1877
rect 1400 2761 1434 2781
rect 1400 2747 1434 2761
rect 1400 2693 1434 2709
rect 1400 2675 1434 2693
rect 1400 2625 1434 2637
rect 1400 2603 1434 2625
rect 1400 2557 1434 2564
rect 1400 2530 1434 2557
rect 1400 2489 1434 2491
rect 1400 2457 1434 2489
rect 1400 2387 1434 2418
rect 1400 2384 1434 2387
rect 1400 2319 1434 2345
rect 1400 2311 1434 2319
rect 1400 2251 1434 2272
rect 1400 2238 1434 2251
rect 1400 2183 1434 2199
rect 1400 2165 1434 2183
rect 1400 2115 1434 2126
rect 1400 2092 1434 2115
rect 1400 2047 1434 2053
rect 1400 2019 1434 2047
rect 1400 1979 1434 1980
rect 1400 1946 1434 1979
rect 1400 1877 1434 1907
rect 1400 1873 1434 1877
rect 1616 2819 1650 2853
rect 1928 2819 1962 2853
rect 1616 2761 1650 2781
rect 1616 2747 1650 2761
rect 1616 2693 1650 2709
rect 1616 2675 1650 2693
rect 1616 2625 1650 2637
rect 1616 2603 1650 2625
rect 1616 2557 1650 2564
rect 1616 2530 1650 2557
rect 1616 2489 1650 2491
rect 1616 2457 1650 2489
rect 1616 2387 1650 2418
rect 1616 2384 1650 2387
rect 1616 2319 1650 2345
rect 1616 2311 1650 2319
rect 1616 2251 1650 2272
rect 1616 2238 1650 2251
rect 1616 2183 1650 2199
rect 1616 2165 1650 2183
rect 1616 2115 1650 2126
rect 1616 2092 1650 2115
rect 1616 2047 1650 2053
rect 1616 2019 1650 2047
rect 1616 1979 1650 1980
rect 1616 1946 1650 1979
rect 1616 1877 1650 1907
rect 1616 1873 1650 1877
rect 1772 2727 1806 2736
rect 1772 2702 1806 2727
rect 1772 2659 1806 2661
rect 1772 2627 1806 2659
rect 1772 2557 1806 2586
rect 1772 2552 1806 2557
rect 1772 2489 1806 2511
rect 1772 2477 1806 2489
rect 1772 2421 1806 2436
rect 1772 2402 1806 2421
rect 1772 2353 1806 2361
rect 1772 2327 1806 2353
rect 1772 2285 1806 2286
rect 1772 2252 1806 2285
rect 1772 2183 1806 2211
rect 1772 2177 1806 2183
rect 1772 2115 1806 2135
rect 1772 2101 1806 2115
rect 1772 2047 1806 2059
rect 1772 2025 1806 2047
rect 1772 1979 1806 1983
rect 1772 1949 1806 1979
rect 1772 1877 1806 1907
rect 1772 1873 1806 1877
rect 2240 2819 2274 2853
rect 1928 2761 1962 2781
rect 1928 2747 1962 2761
rect 1928 2693 1962 2709
rect 1928 2675 1962 2693
rect 1928 2625 1962 2637
rect 1928 2603 1962 2625
rect 1928 2557 1962 2564
rect 1928 2530 1962 2557
rect 1928 2489 1962 2491
rect 1928 2457 1962 2489
rect 1928 2387 1962 2418
rect 1928 2384 1962 2387
rect 1928 2319 1962 2345
rect 1928 2311 1962 2319
rect 1928 2251 1962 2272
rect 1928 2238 1962 2251
rect 1928 2183 1962 2199
rect 1928 2165 1962 2183
rect 1928 2115 1962 2126
rect 1928 2092 1962 2115
rect 1928 2047 1962 2053
rect 1928 2019 1962 2047
rect 1928 1979 1962 1980
rect 1928 1946 1962 1979
rect 1928 1877 1962 1907
rect 1928 1873 1962 1877
rect 2084 2727 2118 2736
rect 2084 2702 2118 2727
rect 2084 2659 2118 2661
rect 2084 2627 2118 2659
rect 2084 2557 2118 2586
rect 2084 2552 2118 2557
rect 2084 2489 2118 2511
rect 2084 2477 2118 2489
rect 2084 2421 2118 2436
rect 2084 2402 2118 2421
rect 2084 2353 2118 2361
rect 2084 2327 2118 2353
rect 2084 2285 2118 2286
rect 2084 2252 2118 2285
rect 2084 2183 2118 2211
rect 2084 2177 2118 2183
rect 2084 2115 2118 2135
rect 2084 2101 2118 2115
rect 2084 2047 2118 2059
rect 2084 2025 2118 2047
rect 2084 1979 2118 1983
rect 2084 1949 2118 1979
rect 2084 1877 2118 1907
rect 2084 1873 2118 1877
rect 2928 2819 2962 2853
rect 2240 2761 2274 2781
rect 2240 2747 2274 2761
rect 2240 2693 2274 2709
rect 2240 2675 2274 2693
rect 2240 2625 2274 2637
rect 2240 2603 2274 2625
rect 2240 2557 2274 2564
rect 2240 2530 2274 2557
rect 2240 2489 2274 2491
rect 2240 2457 2274 2489
rect 2240 2387 2274 2418
rect 2240 2384 2274 2387
rect 2240 2319 2274 2345
rect 2240 2311 2274 2319
rect 2240 2251 2274 2272
rect 2240 2238 2274 2251
rect 2240 2183 2274 2199
rect 2240 2165 2274 2183
rect 2240 2115 2274 2126
rect 2240 2092 2274 2115
rect 2240 2047 2274 2053
rect 2240 2019 2274 2047
rect 2240 1979 2274 1980
rect 2240 1946 2274 1979
rect 2240 1877 2274 1907
rect 2240 1873 2274 1877
rect 2396 2727 2430 2736
rect 2396 2702 2430 2727
rect 2396 2659 2430 2661
rect 2396 2627 2430 2659
rect 2396 2557 2430 2586
rect 2396 2552 2430 2557
rect 2396 2489 2430 2511
rect 2396 2477 2430 2489
rect 2396 2421 2430 2436
rect 2396 2402 2430 2421
rect 2772 2727 2806 2736
rect 2772 2702 2806 2727
rect 2772 2625 2806 2658
rect 2772 2624 2806 2625
rect 2772 2557 2806 2580
rect 2772 2546 2806 2557
rect 2772 2489 2806 2502
rect 2772 2468 2806 2489
rect 2772 2421 2806 2424
rect 2396 2353 2430 2361
rect 2396 2327 2430 2353
rect 2396 2285 2430 2286
rect 2396 2252 2430 2285
rect 2396 2183 2430 2211
rect 2396 2177 2430 2183
rect 2396 2115 2430 2135
rect 2396 2101 2430 2115
rect 2396 2047 2430 2059
rect 2396 2025 2430 2047
rect 2396 1979 2430 1983
rect 2396 1949 2430 1979
rect 2396 1877 2430 1907
rect 2396 1873 2430 1877
rect 2506 2353 2540 2366
rect 2506 2332 2540 2353
rect 2506 2251 2540 2281
rect 2506 2247 2540 2251
rect 2506 2183 2540 2196
rect 2506 2162 2540 2183
rect 2506 2081 2540 2111
rect 2506 2077 2540 2081
rect 2506 2013 2540 2026
rect 2506 1992 2540 2013
rect 2506 1911 2540 1941
rect 2506 1907 2540 1911
rect 2662 2353 2696 2366
rect 2662 2332 2696 2353
rect 2662 2251 2696 2281
rect 2662 2247 2696 2251
rect 2662 2183 2696 2196
rect 2662 2162 2696 2183
rect 2662 2081 2696 2111
rect 2662 2077 2696 2081
rect 2662 2013 2696 2026
rect 2662 1992 2696 2013
rect 2662 1911 2696 1941
rect 2662 1907 2696 1911
rect 2772 2390 2806 2421
rect 2772 2319 2806 2346
rect 2772 2312 2806 2319
rect 2772 2251 2806 2267
rect 2772 2233 2806 2251
rect 2772 2183 2806 2188
rect 2772 2154 2806 2183
rect 2772 2081 2806 2109
rect 2772 2075 2806 2081
rect 2772 2013 2806 2030
rect 2772 1996 2806 2013
rect 2928 2761 2962 2776
rect 2928 2742 2962 2761
rect 2928 2693 2962 2699
rect 2928 2665 2962 2693
rect 2928 2591 2962 2621
rect 2928 2587 2962 2591
rect 2928 2523 2962 2543
rect 2928 2509 2962 2523
rect 2928 2455 2962 2465
rect 2928 2431 2962 2455
rect 2928 2353 2962 2387
rect 2928 2285 2962 2309
rect 2928 2275 2962 2285
rect 2928 2217 2962 2231
rect 2928 2197 2962 2217
rect 2928 2149 2962 2153
rect 2928 2119 2962 2149
rect 2928 2047 2962 2075
rect 2928 2041 2962 2047
rect 2928 1979 2962 1997
rect 2928 1963 2962 1979
rect 3084 2727 3118 2736
rect 3084 2702 3118 2727
rect 3084 2659 3118 2661
rect 3084 2627 3118 2659
rect 3084 2557 3118 2586
rect 3084 2552 3118 2557
rect 3084 2489 3118 2511
rect 3084 2477 3118 2489
rect 3084 2421 3118 2436
rect 3084 2402 3118 2421
rect 3458 2405 3492 2439
rect 3530 2405 3564 2439
rect 3084 2353 3118 2361
rect 3084 2327 3118 2353
rect 3646 2325 3680 2359
rect 3084 2285 3118 2286
rect 3084 2252 3118 2285
rect 3396 2262 3430 2296
rect 3468 2262 3502 2296
rect 3646 2253 3680 2287
rect 3791 2337 3825 2371
rect 3791 2265 3825 2299
rect 3894 2324 3928 2358
rect 3894 2252 3928 2286
rect 3084 2183 3118 2211
rect 3084 2177 3118 2183
rect 3084 2115 3118 2136
rect 3084 2102 3118 2115
rect 3084 2047 3118 2060
rect 3084 2026 3118 2047
rect 3084 1979 3118 1984
rect 3084 1950 3118 1979
rect 137 1783 169 1817
rect 169 1783 171 1817
rect 231 1783 264 1817
rect 264 1783 265 1817
rect 324 1783 325 1817
rect 325 1783 358 1817
rect 578 1783 591 1817
rect 591 1783 612 1817
rect 650 1783 651 1817
rect 651 1783 684 1817
rect 784 1783 807 1817
rect 807 1783 818 1817
rect 856 1783 867 1817
rect 867 1783 890 1817
rect 985 1783 989 1817
rect 989 1783 1019 1817
rect 1084 1783 1118 1817
rect 1183 1783 1213 1817
rect 1213 1783 1217 1817
rect 1407 1783 1441 1817
rect 1479 1783 1487 1817
rect 1487 1783 1513 1817
rect 1673 1783 1677 1817
rect 1677 1783 1707 1817
rect 1767 1783 1772 1817
rect 1772 1783 1801 1817
rect 1860 1783 1867 1817
rect 1867 1783 1894 1817
rect 1992 1783 2023 1817
rect 2023 1783 2026 1817
rect 2086 1783 2118 1817
rect 2118 1783 2120 1817
rect 2179 1783 2213 1817
rect 2306 1783 2335 1817
rect 2335 1783 2340 1817
rect 2378 1783 2403 1817
rect 2403 1783 2412 1817
rect 2510 1783 2533 1817
rect 2533 1783 2544 1817
rect 2582 1783 2601 1817
rect 2601 1783 2616 1817
rect 2795 1783 2799 1817
rect 2799 1783 2829 1817
rect 2867 1783 2901 1817
rect 2987 1783 2989 1817
rect 2989 1783 3021 1817
rect 3059 1783 3091 1817
rect 3091 1783 3093 1817
rect 112 246 139 280
rect 139 246 146 280
rect 189 246 208 280
rect 208 246 223 280
rect 266 246 277 280
rect 277 246 300 280
rect 343 246 346 280
rect 346 246 377 280
rect 420 246 450 280
rect 450 246 454 280
rect 497 246 519 280
rect 519 246 531 280
rect 574 246 587 280
rect 587 246 608 280
rect 651 246 655 280
rect 655 246 685 280
rect 728 246 757 280
rect 757 246 762 280
rect 805 246 825 280
rect 825 246 839 280
rect 882 246 893 280
rect 893 246 916 280
rect 958 246 961 280
rect 961 246 992 280
rect 1034 246 1063 280
rect 1063 246 1068 280
rect 1198 246 1219 280
rect 1219 246 1232 280
rect 1270 246 1279 280
rect 1279 246 1304 280
rect 1415 246 1435 280
rect 1435 246 1449 280
rect 1492 246 1504 280
rect 1504 246 1526 280
rect 1569 246 1573 280
rect 1573 246 1603 280
rect 1646 246 1677 280
rect 1677 246 1680 280
rect 1723 246 1746 280
rect 1746 246 1757 280
rect 1800 246 1815 280
rect 1815 246 1834 280
rect 1877 246 1883 280
rect 1883 246 1911 280
rect 1954 246 1985 280
rect 1985 246 1988 280
rect 2031 246 2053 280
rect 2053 246 2065 280
rect 2108 246 2121 280
rect 2121 246 2142 280
rect 2185 246 2189 280
rect 2189 246 2219 280
rect 2261 246 2291 280
rect 2291 246 2295 280
rect 2337 246 2359 280
rect 2359 246 2371 280
rect 2507 246 2515 280
rect 2515 246 2541 280
rect 2585 246 2590 280
rect 2590 246 2619 280
rect 2663 246 2665 280
rect 2665 246 2697 280
rect 2741 246 2775 280
rect 2819 246 2853 280
rect 2896 246 2927 280
rect 2927 246 2930 280
rect 2973 246 3001 280
rect 3001 246 3007 280
rect 3050 246 3075 280
rect 3075 246 3084 280
rect 3127 246 3149 280
rect 3149 246 3161 280
rect 3204 246 3223 280
rect 3223 246 3238 280
rect 3473 246 3489 280
rect 3489 246 3507 280
rect 3545 246 3549 280
rect 3549 246 3579 280
rect 3799 246 3815 280
rect 3815 246 3833 280
rect 3871 246 3875 280
rect 3875 246 3905 280
rect 4125 246 4141 280
rect 4141 246 4159 280
rect 4197 246 4201 280
rect 4201 246 4231 280
rect 4489 258 4508 285
rect 4508 258 4523 285
rect 4562 258 4583 285
rect 4583 258 4596 285
rect 4635 258 4657 285
rect 4657 258 4669 285
rect 4708 258 4731 285
rect 4731 258 4742 285
rect 4781 258 4805 285
rect 4805 258 4815 285
rect 4854 258 4879 285
rect 4879 258 4888 285
rect 4926 258 4953 285
rect 4953 258 4960 285
rect 4998 258 5027 285
rect 5027 258 5032 285
rect 5070 258 5101 285
rect 5101 258 5104 285
rect 5142 258 5175 285
rect 5175 258 5176 285
rect 4489 251 4523 258
rect 4562 251 4596 258
rect 4635 251 4669 258
rect 4708 251 4742 258
rect 4781 251 4815 258
rect 4854 251 4888 258
rect 4926 251 4960 258
rect 4998 251 5032 258
rect 5070 251 5104 258
rect 5142 251 5176 258
rect 5360 246 5389 280
rect 5389 246 5394 280
rect 5433 246 5457 280
rect 5457 246 5467 280
rect 5577 246 5579 280
rect 5579 246 5611 280
rect 5649 246 5681 280
rect 5681 246 5683 280
rect 44 162 78 196
rect 44 94 78 122
rect 44 88 78 94
rect 44 26 78 48
rect 44 14 78 26
rect 44 -42 78 -26
rect 44 -60 78 -42
rect 44 -110 78 -100
rect 44 -134 78 -110
rect 44 -178 78 -174
rect 44 -208 78 -178
rect 44 -280 78 -248
rect 44 -282 78 -280
rect 44 -348 78 -322
rect 44 -356 78 -348
rect 44 -416 78 -395
rect 44 -429 78 -416
rect 44 -484 78 -468
rect 44 -502 78 -484
rect 44 -552 78 -541
rect 44 -575 78 -552
rect 44 -620 78 -614
rect 44 -648 78 -620
rect 44 -688 78 -687
rect 44 -721 78 -688
rect 44 -790 78 -760
rect 44 -794 78 -790
rect 260 162 294 196
rect 692 162 726 196
rect 260 94 294 121
rect 260 87 294 94
rect 260 26 294 46
rect 260 12 294 26
rect 260 -42 294 -29
rect 260 -63 294 -42
rect 260 -110 294 -104
rect 260 -138 294 -110
rect 260 -212 294 -179
rect 260 -213 294 -212
rect 260 -280 294 -254
rect 260 -288 294 -280
rect 260 -348 294 -329
rect 260 -363 294 -348
rect 260 -416 294 -404
rect 260 -438 294 -416
rect 260 -484 294 -479
rect 260 -513 294 -484
rect 260 -586 294 -554
rect 260 -588 294 -586
rect 260 -654 294 -628
rect 260 -662 294 -654
rect 476 60 510 64
rect 476 30 510 60
rect 476 -42 510 -11
rect 476 -45 510 -42
rect 476 -110 510 -86
rect 476 -120 510 -110
rect 476 -178 510 -161
rect 476 -195 510 -178
rect 476 -246 510 -236
rect 476 -270 510 -246
rect 476 -314 510 -311
rect 476 -345 510 -314
rect 476 -416 510 -386
rect 476 -420 510 -416
rect 476 -484 510 -461
rect 476 -495 510 -484
rect 476 -552 510 -536
rect 476 -570 510 -552
rect 476 -620 510 -611
rect 476 -645 510 -620
rect 476 -688 510 -686
rect 476 -720 510 -688
rect 476 -790 510 -760
rect 476 -794 510 -790
rect 1124 162 1158 196
rect 692 94 726 121
rect 692 87 726 94
rect 692 26 726 46
rect 692 12 726 26
rect 692 -42 726 -29
rect 692 -63 726 -42
rect 692 -110 726 -104
rect 692 -138 726 -110
rect 692 -212 726 -179
rect 692 -213 726 -212
rect 692 -280 726 -254
rect 692 -288 726 -280
rect 692 -348 726 -329
rect 692 -363 726 -348
rect 692 -416 726 -404
rect 692 -438 726 -416
rect 692 -484 726 -479
rect 692 -513 726 -484
rect 692 -586 726 -554
rect 692 -588 726 -586
rect 692 -654 726 -628
rect 692 -662 726 -654
rect 908 60 942 64
rect 908 30 942 60
rect 908 -42 942 -11
rect 908 -45 942 -42
rect 908 -110 942 -86
rect 908 -120 942 -110
rect 908 -178 942 -161
rect 908 -195 942 -178
rect 908 -246 942 -236
rect 908 -270 942 -246
rect 908 -314 942 -311
rect 908 -345 942 -314
rect 908 -416 942 -386
rect 908 -420 942 -416
rect 908 -484 942 -461
rect 908 -495 942 -484
rect 908 -552 942 -536
rect 908 -570 942 -552
rect 908 -620 942 -611
rect 908 -645 942 -620
rect 908 -688 942 -686
rect 908 -720 942 -688
rect 908 -790 942 -760
rect 908 -794 942 -790
rect 1556 162 1590 196
rect 1124 94 1158 121
rect 1124 87 1158 94
rect 1124 26 1158 46
rect 1124 12 1158 26
rect 1124 -42 1158 -29
rect 1124 -63 1158 -42
rect 1124 -110 1158 -104
rect 1124 -138 1158 -110
rect 1124 -212 1158 -179
rect 1124 -213 1158 -212
rect 1124 -280 1158 -254
rect 1124 -288 1158 -280
rect 1124 -348 1158 -329
rect 1124 -363 1158 -348
rect 1124 -416 1158 -404
rect 1124 -438 1158 -416
rect 1124 -484 1158 -479
rect 1124 -513 1158 -484
rect 1124 -586 1158 -554
rect 1124 -588 1158 -586
rect 1124 -654 1158 -628
rect 1124 -662 1158 -654
rect 1340 60 1374 64
rect 1340 30 1374 60
rect 1340 -42 1374 -11
rect 1340 -45 1374 -42
rect 1340 -110 1374 -86
rect 1340 -120 1374 -110
rect 1340 -178 1374 -161
rect 1340 -195 1374 -178
rect 1340 -246 1374 -236
rect 1340 -270 1374 -246
rect 1340 -314 1374 -311
rect 1340 -345 1374 -314
rect 1340 -416 1374 -386
rect 1340 -420 1374 -416
rect 1340 -484 1374 -461
rect 1340 -495 1374 -484
rect 1340 -552 1374 -536
rect 1340 -570 1374 -552
rect 1340 -620 1374 -611
rect 1340 -645 1374 -620
rect 1340 -688 1374 -686
rect 1340 -720 1374 -688
rect 1340 -790 1374 -760
rect 1340 -794 1374 -790
rect 1988 162 2022 196
rect 1556 94 1590 121
rect 1556 87 1590 94
rect 1556 26 1590 46
rect 1556 12 1590 26
rect 1556 -42 1590 -29
rect 1556 -63 1590 -42
rect 1556 -110 1590 -104
rect 1556 -138 1590 -110
rect 1556 -212 1590 -179
rect 1556 -213 1590 -212
rect 1556 -280 1590 -254
rect 1556 -288 1590 -280
rect 1556 -348 1590 -329
rect 1556 -363 1590 -348
rect 1556 -416 1590 -404
rect 1556 -438 1590 -416
rect 1556 -484 1590 -479
rect 1556 -513 1590 -484
rect 1556 -586 1590 -554
rect 1556 -588 1590 -586
rect 1556 -654 1590 -628
rect 1556 -662 1590 -654
rect 1772 60 1806 64
rect 1772 30 1806 60
rect 1772 -42 1806 -11
rect 1772 -45 1806 -42
rect 1772 -110 1806 -86
rect 1772 -120 1806 -110
rect 1772 -178 1806 -161
rect 1772 -195 1806 -178
rect 1772 -246 1806 -236
rect 1772 -270 1806 -246
rect 1772 -314 1806 -311
rect 1772 -345 1806 -314
rect 1772 -416 1806 -386
rect 1772 -420 1806 -416
rect 1772 -484 1806 -461
rect 1772 -495 1806 -484
rect 1772 -552 1806 -536
rect 1772 -570 1806 -552
rect 1772 -620 1806 -611
rect 1772 -645 1806 -620
rect 1772 -688 1806 -686
rect 1772 -720 1806 -688
rect 1772 -790 1806 -760
rect 1772 -794 1806 -790
rect 2420 162 2454 196
rect 1988 94 2022 121
rect 1988 87 2022 94
rect 1988 26 2022 46
rect 1988 12 2022 26
rect 1988 -42 2022 -29
rect 1988 -63 2022 -42
rect 1988 -110 2022 -104
rect 1988 -138 2022 -110
rect 1988 -212 2022 -179
rect 1988 -213 2022 -212
rect 1988 -280 2022 -254
rect 1988 -288 2022 -280
rect 1988 -348 2022 -329
rect 1988 -363 2022 -348
rect 1988 -416 2022 -404
rect 1988 -438 2022 -416
rect 1988 -484 2022 -479
rect 1988 -513 2022 -484
rect 1988 -586 2022 -554
rect 1988 -588 2022 -586
rect 1988 -654 2022 -628
rect 1988 -662 2022 -654
rect 2204 60 2238 64
rect 2204 30 2238 60
rect 2204 -42 2238 -11
rect 2204 -45 2238 -42
rect 2204 -110 2238 -86
rect 2204 -120 2238 -110
rect 2204 -178 2238 -161
rect 2204 -195 2238 -178
rect 2204 -246 2238 -236
rect 2204 -270 2238 -246
rect 2204 -314 2238 -311
rect 2204 -345 2238 -314
rect 2204 -416 2238 -386
rect 2204 -420 2238 -416
rect 2204 -484 2238 -461
rect 2204 -495 2238 -484
rect 2204 -552 2238 -536
rect 2204 -570 2238 -552
rect 2204 -620 2238 -611
rect 2204 -645 2238 -620
rect 2204 -688 2238 -686
rect 2204 -720 2238 -688
rect 2204 -790 2238 -760
rect 2204 -794 2238 -790
rect 2852 162 2886 196
rect 2420 94 2454 121
rect 2420 87 2454 94
rect 2420 26 2454 46
rect 2420 12 2454 26
rect 2420 -42 2454 -29
rect 2420 -63 2454 -42
rect 2420 -110 2454 -104
rect 2420 -138 2454 -110
rect 2420 -212 2454 -179
rect 2420 -213 2454 -212
rect 2420 -280 2454 -254
rect 2420 -288 2454 -280
rect 2420 -348 2454 -329
rect 2420 -363 2454 -348
rect 2420 -416 2454 -404
rect 2420 -438 2454 -416
rect 2420 -484 2454 -479
rect 2420 -513 2454 -484
rect 2420 -586 2454 -554
rect 2420 -588 2454 -586
rect 2420 -654 2454 -628
rect 2420 -662 2454 -654
rect 2636 60 2670 64
rect 2636 30 2670 60
rect 2636 -42 2670 -11
rect 2636 -45 2670 -42
rect 2636 -110 2670 -86
rect 2636 -120 2670 -110
rect 2636 -178 2670 -161
rect 2636 -195 2670 -178
rect 2636 -246 2670 -236
rect 2636 -270 2670 -246
rect 2636 -314 2670 -311
rect 2636 -345 2670 -314
rect 2636 -416 2670 -386
rect 2636 -420 2670 -416
rect 2636 -484 2670 -461
rect 2636 -495 2670 -484
rect 2636 -552 2670 -536
rect 2636 -570 2670 -552
rect 2636 -620 2670 -611
rect 2636 -645 2670 -620
rect 2636 -688 2670 -686
rect 2636 -720 2670 -688
rect 2636 -790 2670 -760
rect 2636 -794 2670 -790
rect 3284 162 3318 196
rect 2852 94 2886 121
rect 2852 87 2886 94
rect 2852 26 2886 46
rect 2852 12 2886 26
rect 2852 -42 2886 -29
rect 2852 -63 2886 -42
rect 2852 -110 2886 -104
rect 2852 -138 2886 -110
rect 2852 -212 2886 -179
rect 2852 -213 2886 -212
rect 2852 -280 2886 -254
rect 2852 -288 2886 -280
rect 2852 -348 2886 -329
rect 2852 -363 2886 -348
rect 2852 -416 2886 -404
rect 2852 -438 2886 -416
rect 2852 -484 2886 -479
rect 2852 -513 2886 -484
rect 2852 -586 2886 -554
rect 2852 -588 2886 -586
rect 2852 -654 2886 -628
rect 2852 -662 2886 -654
rect 3068 60 3102 64
rect 3068 30 3102 60
rect 3068 -42 3102 -11
rect 3068 -45 3102 -42
rect 3068 -110 3102 -86
rect 3068 -120 3102 -110
rect 3068 -178 3102 -161
rect 3068 -195 3102 -178
rect 3068 -246 3102 -236
rect 3068 -270 3102 -246
rect 3068 -314 3102 -311
rect 3068 -345 3102 -314
rect 3068 -416 3102 -386
rect 3068 -420 3102 -416
rect 3068 -484 3102 -461
rect 3068 -495 3102 -484
rect 3068 -552 3102 -536
rect 3068 -570 3102 -552
rect 3068 -620 3102 -611
rect 3068 -645 3102 -620
rect 3068 -688 3102 -686
rect 3068 -720 3102 -688
rect 3068 -790 3102 -760
rect 3068 -794 3102 -790
rect 3284 94 3318 121
rect 3284 87 3318 94
rect 3284 26 3318 46
rect 3284 12 3318 26
rect 3284 -42 3318 -29
rect 3284 -63 3318 -42
rect 3284 -110 3318 -104
rect 3284 -138 3318 -110
rect 3284 -212 3318 -179
rect 3284 -213 3318 -212
rect 3284 -280 3318 -254
rect 3284 -288 3318 -280
rect 3284 -348 3318 -329
rect 3284 -363 3318 -348
rect 3284 -416 3318 -404
rect 3284 -438 3318 -416
rect 3284 -484 3318 -479
rect 3284 -513 3318 -484
rect 3284 -586 3318 -554
rect 3284 -588 3318 -586
rect 3284 -654 3318 -628
rect 3284 -662 3318 -654
rect 3394 162 3428 196
rect 4372 167 4406 196
rect 4372 162 4406 167
rect 3394 94 3428 121
rect 3394 87 3428 94
rect 3394 26 3428 46
rect 3394 12 3428 26
rect 3394 -42 3428 -29
rect 3394 -63 3428 -42
rect 3394 -110 3428 -104
rect 3394 -138 3428 -110
rect 3394 -212 3428 -179
rect 3394 -213 3428 -212
rect 3394 -280 3428 -254
rect 3394 -288 3428 -280
rect 3394 -348 3428 -329
rect 3394 -363 3428 -348
rect 3394 -416 3428 -404
rect 3394 -438 3428 -416
rect 3394 -484 3428 -479
rect 3394 -513 3428 -484
rect 3394 -586 3428 -554
rect 3394 -588 3428 -586
rect 3394 -654 3428 -628
rect 3394 -662 3428 -654
rect 3610 60 3644 64
rect 3610 30 3644 60
rect 3610 -42 3644 -11
rect 3610 -45 3644 -42
rect 3610 -110 3644 -86
rect 3610 -120 3644 -110
rect 3610 -178 3644 -161
rect 3610 -195 3644 -178
rect 3610 -246 3644 -236
rect 3610 -270 3644 -246
rect 3610 -314 3644 -311
rect 3610 -345 3644 -314
rect 3610 -416 3644 -386
rect 3610 -420 3644 -416
rect 3610 -484 3644 -461
rect 3610 -495 3644 -484
rect 3610 -552 3644 -536
rect 3610 -570 3644 -552
rect 3610 -620 3644 -611
rect 3610 -645 3644 -620
rect 3610 -688 3644 -686
rect 3610 -720 3644 -688
rect 3610 -790 3644 -760
rect 3610 -794 3644 -790
rect 3720 60 3754 64
rect 3720 30 3754 60
rect 3720 -42 3754 -11
rect 3720 -45 3754 -42
rect 3720 -110 3754 -86
rect 3720 -120 3754 -110
rect 3720 -178 3754 -161
rect 3720 -195 3754 -178
rect 3720 -246 3754 -236
rect 3720 -270 3754 -246
rect 3720 -314 3754 -311
rect 3720 -345 3754 -314
rect 3720 -416 3754 -386
rect 3720 -420 3754 -416
rect 3720 -484 3754 -461
rect 3720 -495 3754 -484
rect 3720 -552 3754 -536
rect 3720 -570 3754 -552
rect 3720 -620 3754 -611
rect 3720 -645 3754 -620
rect 3720 -688 3754 -686
rect 3720 -720 3754 -688
rect 3720 -790 3754 -760
rect 3720 -794 3754 -790
rect 3936 60 3970 64
rect 3936 30 3970 60
rect 3936 -42 3970 -11
rect 3936 -45 3970 -42
rect 3936 -110 3970 -86
rect 3936 -120 3970 -110
rect 3936 -178 3970 -161
rect 3936 -195 3970 -178
rect 3936 -246 3970 -236
rect 3936 -270 3970 -246
rect 3936 -314 3970 -311
rect 3936 -345 3970 -314
rect 3936 -416 3970 -386
rect 3936 -420 3970 -416
rect 3936 -484 3970 -461
rect 3936 -495 3970 -484
rect 3936 -552 3970 -536
rect 3936 -570 3970 -552
rect 3936 -620 3970 -611
rect 3936 -645 3970 -620
rect 3936 -688 3970 -686
rect 3936 -720 3970 -688
rect 3936 -790 3970 -760
rect 3936 -794 3970 -790
rect 4046 60 4080 64
rect 4046 30 4080 60
rect 4046 -42 4080 -11
rect 4046 -45 4080 -42
rect 4046 -110 4080 -86
rect 4046 -120 4080 -110
rect 4046 -178 4080 -161
rect 4046 -195 4080 -178
rect 4046 -246 4080 -236
rect 4046 -270 4080 -246
rect 4046 -314 4080 -311
rect 4046 -345 4080 -314
rect 4046 -416 4080 -386
rect 4046 -420 4080 -416
rect 4046 -484 4080 -461
rect 4046 -495 4080 -484
rect 4046 -552 4080 -536
rect 4046 -570 4080 -552
rect 4046 -620 4080 -611
rect 4046 -645 4080 -620
rect 4046 -688 4080 -686
rect 4046 -720 4080 -688
rect 4046 -790 4080 -760
rect 4046 -794 4080 -790
rect 4262 60 4296 64
rect 4262 30 4296 60
rect 4372 99 4406 124
rect 4372 90 4406 99
rect 4552 7 4586 41
rect 4804 167 4838 196
rect 4804 162 4838 167
rect 4804 99 4838 124
rect 4804 90 4838 99
rect 4624 7 4658 41
rect 4984 7 5018 41
rect 5236 167 5270 196
rect 5236 162 5270 167
rect 5236 99 5270 124
rect 5236 90 5270 99
rect 5056 7 5090 41
rect 4262 -42 4296 -11
rect 4262 -45 4296 -42
rect 4262 -110 4296 -86
rect 4262 -120 4296 -110
rect 5362 -8 5396 19
rect 5362 -15 5396 -8
rect 5362 -76 5396 -56
rect 5362 -90 5396 -76
rect 4685 -120 4719 -119
rect 4777 -120 4811 -119
rect 4868 -120 4902 -119
rect 4471 -154 4505 -120
rect 4543 -154 4567 -120
rect 4567 -154 4577 -120
rect 4685 -153 4689 -120
rect 4689 -153 4719 -120
rect 4777 -153 4784 -120
rect 4784 -153 4811 -120
rect 4868 -153 4879 -120
rect 4879 -153 4902 -120
rect 4997 -154 5001 -120
rect 5001 -154 5031 -120
rect 5081 -154 5096 -120
rect 5096 -154 5115 -120
rect 5165 -154 5191 -120
rect 5191 -154 5199 -120
rect 5362 -144 5396 -131
rect 4262 -178 4296 -161
rect 4262 -195 4296 -178
rect 4262 -246 4296 -236
rect 4262 -270 4296 -246
rect 5362 -165 5396 -144
rect 5362 -212 5396 -206
rect 5362 -240 5396 -212
rect 4262 -314 4296 -311
rect 4262 -345 4296 -314
rect 4262 -416 4296 -386
rect 4262 -420 4296 -416
rect 4262 -484 4296 -461
rect 4262 -495 4296 -484
rect 4262 -552 4296 -536
rect 4262 -570 4296 -552
rect 4262 -620 4296 -611
rect 4262 -645 4296 -620
rect 4262 -688 4296 -686
rect 4262 -720 4296 -688
rect 4262 -790 4296 -760
rect 4262 -794 4296 -790
rect 4372 -280 4406 -264
rect 4372 -298 4406 -280
rect 4372 -348 4406 -339
rect 4372 -373 4406 -348
rect 4372 -416 4406 -415
rect 4372 -449 4406 -416
rect 4372 -518 4406 -491
rect 4372 -525 4406 -518
rect 4372 -586 4406 -567
rect 4372 -601 4406 -586
rect 4372 -654 4406 -643
rect 4372 -677 4406 -654
rect 4628 -382 4662 -381
rect 4628 -415 4662 -382
rect 4628 -484 4662 -456
rect 4628 -490 4662 -484
rect 4628 -552 4662 -532
rect 4628 -566 4662 -552
rect 4628 -620 4662 -608
rect 4628 -642 4662 -620
rect 4628 -688 4662 -684
rect 4628 -718 4662 -688
rect 4628 -790 4662 -760
rect 4628 -794 4662 -790
rect 4784 -280 4818 -276
rect 4784 -310 4818 -280
rect 4784 -382 4818 -351
rect 4784 -385 4818 -382
rect 4784 -450 4818 -427
rect 4784 -461 4818 -450
rect 4784 -518 4818 -503
rect 4784 -537 4818 -518
rect 4784 -586 4818 -579
rect 4784 -613 4818 -586
rect 4784 -688 4818 -655
rect 4784 -689 4818 -688
rect 4940 -382 4974 -381
rect 4940 -415 4974 -382
rect 4940 -484 4974 -456
rect 4940 -490 4974 -484
rect 4940 -552 4974 -532
rect 4940 -566 4974 -552
rect 4940 -620 4974 -608
rect 4940 -642 4974 -620
rect 4940 -688 4974 -684
rect 4940 -718 4974 -688
rect 4940 -790 4974 -760
rect 4940 -794 4974 -790
rect 5096 -280 5130 -276
rect 5096 -310 5130 -280
rect 5096 -382 5130 -351
rect 5096 -385 5130 -382
rect 5096 -450 5130 -427
rect 5096 -461 5130 -450
rect 5096 -518 5130 -503
rect 5096 -537 5130 -518
rect 5096 -586 5130 -579
rect 5096 -613 5130 -586
rect 5096 -688 5130 -655
rect 5096 -689 5130 -688
rect 5252 -382 5286 -381
rect 5252 -415 5286 -382
rect 5252 -484 5286 -456
rect 5252 -490 5286 -484
rect 5252 -552 5286 -532
rect 5252 -566 5286 -552
rect 5252 -620 5286 -608
rect 5252 -642 5286 -620
rect 5252 -688 5286 -684
rect 5252 -718 5286 -688
rect 5252 -790 5286 -760
rect 5252 -794 5286 -790
rect 5362 -314 5396 -281
rect 5362 -315 5396 -314
rect 5362 -382 5396 -356
rect 5362 -390 5396 -382
rect 5362 -450 5396 -431
rect 5362 -465 5396 -450
rect 5362 -518 5396 -506
rect 5362 -540 5396 -518
rect 5362 -586 5396 -582
rect 5362 -616 5396 -586
rect 5518 -8 5552 19
rect 5518 -15 5552 -8
rect 5518 -76 5552 -58
rect 5518 -92 5552 -76
rect 5518 -144 5552 -136
rect 5518 -170 5552 -144
rect 5518 -246 5552 -214
rect 5518 -248 5552 -246
rect 5518 -314 5552 -292
rect 5518 -326 5552 -314
rect 5518 -382 5552 -370
rect 5518 -404 5552 -382
rect 5518 -450 5552 -448
rect 5518 -482 5552 -450
rect 5518 -552 5552 -526
rect 5518 -560 5552 -552
rect 5518 -620 5552 -604
rect 5518 -638 5552 -620
rect 5518 -688 5552 -682
rect 5518 -716 5552 -688
rect 5518 -790 5552 -760
rect 5518 -794 5552 -790
rect 5675 94 5708 109
rect 5708 94 5709 109
rect 5675 75 5709 94
rect 5675 26 5708 33
rect 5708 26 5709 33
rect 5675 -1 5709 26
rect 5675 -76 5709 -43
rect 5675 -77 5708 -76
rect 5708 -77 5709 -76
rect 5675 -144 5709 -120
rect 5675 -154 5708 -144
rect 5708 -154 5709 -144
rect 5675 -212 5709 -197
rect 5675 -231 5708 -212
rect 5708 -231 5709 -212
rect 5675 -280 5709 -274
rect 5675 -308 5708 -280
rect 5708 -308 5709 -280
rect 5675 -382 5708 -351
rect 5708 -382 5709 -351
rect 5675 -385 5709 -382
rect 5675 -450 5708 -428
rect 5708 -450 5709 -428
rect 5675 -462 5709 -450
rect 5675 -518 5708 -505
rect 5708 -518 5709 -505
rect 5675 -539 5709 -518
rect 5675 -586 5708 -582
rect 5708 -586 5709 -582
rect 5675 -616 5709 -586
rect 67 -912 91 -878
rect 91 -912 101 -878
rect 140 -912 160 -878
rect 160 -912 174 -878
rect 213 -912 229 -878
rect 229 -912 247 -878
rect 286 -912 298 -878
rect 298 -912 320 -878
rect 359 -912 367 -878
rect 367 -912 393 -878
rect 432 -912 436 -878
rect 436 -912 466 -878
rect 505 -912 539 -878
rect 578 -912 608 -878
rect 608 -912 612 -878
rect 651 -912 677 -878
rect 677 -912 685 -878
rect 724 -912 746 -878
rect 746 -912 758 -878
rect 797 -912 815 -878
rect 815 -912 831 -878
rect 870 -912 884 -878
rect 884 -912 904 -878
rect 943 -912 953 -878
rect 953 -912 977 -878
rect 1016 -912 1022 -878
rect 1022 -912 1050 -878
rect 1089 -912 1091 -878
rect 1091 -912 1123 -878
rect 1162 -912 1195 -878
rect 1195 -912 1196 -878
rect 1235 -912 1264 -878
rect 1264 -912 1269 -878
rect 1308 -912 1333 -878
rect 1333 -912 1342 -878
rect 1381 -912 1402 -878
rect 1402 -912 1415 -878
rect 1454 -912 1471 -878
rect 1471 -912 1488 -878
rect 1527 -912 1540 -878
rect 1540 -912 1561 -878
rect 1600 -912 1609 -878
rect 1609 -912 1634 -878
rect 1673 -912 1678 -878
rect 1678 -912 1707 -878
rect 1746 -912 1747 -878
rect 1747 -912 1780 -878
rect 1819 -912 1850 -878
rect 1850 -912 1853 -878
rect 1892 -912 1919 -878
rect 1919 -912 1926 -878
rect 1965 -912 1988 -878
rect 1988 -912 1999 -878
rect 2038 -912 2057 -878
rect 2057 -912 2072 -878
rect 2111 -912 2126 -878
rect 2126 -912 2145 -878
rect 2184 -912 2195 -878
rect 2195 -912 2218 -878
rect 2257 -912 2264 -878
rect 2264 -912 2291 -878
rect 2330 -912 2333 -878
rect 2333 -912 2364 -878
rect 2403 -912 2437 -878
rect 2476 -912 2505 -878
rect 2505 -912 2510 -878
rect 2549 -912 2573 -878
rect 2573 -912 2583 -878
rect 2622 -912 2641 -878
rect 2641 -912 2656 -878
rect 2695 -912 2709 -878
rect 2709 -912 2729 -878
rect 2768 -912 2777 -878
rect 2777 -912 2802 -878
rect 2841 -912 2845 -878
rect 2845 -912 2875 -878
rect 2914 -912 2947 -878
rect 2947 -912 2948 -878
rect 2987 -912 3015 -878
rect 3015 -912 3021 -878
rect 3060 -912 3083 -878
rect 3083 -912 3094 -878
rect 3133 -912 3151 -878
rect 3151 -912 3167 -878
rect 3206 -912 3219 -878
rect 3219 -912 3240 -878
rect 3279 -912 3287 -878
rect 3287 -912 3313 -878
rect 3352 -912 3355 -878
rect 3355 -912 3386 -878
rect 3425 -912 3457 -878
rect 3457 -912 3459 -878
rect 3498 -912 3525 -878
rect 3525 -912 3532 -878
rect 3570 -912 3593 -878
rect 3593 -912 3604 -878
rect 3642 -912 3661 -878
rect 3661 -912 3676 -878
rect 3714 -912 3729 -878
rect 3729 -912 3748 -878
rect 3786 -912 3797 -878
rect 3797 -912 3820 -878
rect 3858 -912 3865 -878
rect 3865 -912 3892 -878
rect 3930 -912 3933 -878
rect 3933 -912 3964 -878
rect 4002 -912 4035 -878
rect 4035 -912 4036 -878
rect 4074 -912 4103 -878
rect 4103 -912 4108 -878
rect 4146 -912 4171 -878
rect 4171 -912 4180 -878
rect 4218 -912 4239 -878
rect 4239 -912 4252 -878
rect 4290 -912 4307 -878
rect 4307 -912 4324 -878
rect 4362 -912 4375 -878
rect 4375 -912 4396 -878
rect 4434 -912 4443 -878
rect 4443 -912 4468 -878
rect 4506 -912 4511 -878
rect 4511 -912 4540 -878
rect 4578 -912 4579 -878
rect 4579 -912 4612 -878
rect 4650 -912 4681 -878
rect 4681 -912 4684 -878
rect 4722 -912 4749 -878
rect 4749 -912 4756 -878
rect 4794 -912 4817 -878
rect 4817 -912 4828 -878
rect 4866 -912 4885 -878
rect 4885 -912 4900 -878
rect 4938 -912 4953 -878
rect 4953 -912 4972 -878
rect 5010 -912 5021 -878
rect 5021 -912 5044 -878
rect 5082 -912 5089 -878
rect 5089 -912 5116 -878
rect 5154 -912 5157 -878
rect 5157 -912 5188 -878
rect 5226 -912 5259 -878
rect 5259 -912 5260 -878
rect 5298 -912 5327 -878
rect 5327 -912 5332 -878
rect 5370 -912 5395 -878
rect 5395 -912 5404 -878
rect 5442 -912 5463 -878
rect 5463 -912 5476 -878
rect 5514 -912 5531 -878
rect 5531 -912 5548 -878
rect 5586 -912 5599 -878
rect 5599 -912 5620 -878
rect 5658 -912 5667 -878
rect 5667 -912 5692 -878
<< metal1 >>
rect 68 2981 3983 3016
rect 68 2947 80 2981
rect 114 2947 153 2981
rect 187 2947 226 2981
rect 260 2947 299 2981
rect 333 2947 372 2981
rect 406 2947 445 2981
rect 479 2947 518 2981
rect 552 2947 591 2981
rect 625 2947 664 2981
rect 698 2947 737 2981
rect 771 2947 810 2981
rect 844 2947 883 2981
rect 917 2947 956 2981
rect 990 2947 1029 2981
rect 1063 2947 1102 2981
rect 1136 2947 1175 2981
rect 1209 2947 1248 2981
rect 1282 2947 1321 2981
rect 1355 2947 1394 2981
rect 1428 2947 1467 2981
rect 1501 2947 1540 2981
rect 1574 2947 1613 2981
rect 1647 2947 1686 2981
rect 1720 2947 1759 2981
rect 1793 2947 1832 2981
rect 1866 2947 1905 2981
rect 1939 2947 1978 2981
rect 2012 2947 2051 2981
rect 2085 2947 2124 2981
rect 2158 2947 2197 2981
rect 2231 2947 2270 2981
rect 2304 2947 2343 2981
rect 2377 2947 2416 2981
rect 2450 2947 2489 2981
rect 2523 2947 2562 2981
rect 2596 2947 2635 2981
rect 2669 2947 2708 2981
rect 2742 2947 2781 2981
rect 2815 2947 2854 2981
rect 2888 2947 2927 2981
rect 2961 2947 3000 2981
rect 3034 2947 3072 2981
rect 3106 2947 3144 2981
rect 3178 2947 3216 2981
rect 3250 2947 3288 2981
rect 3322 2947 3360 2981
rect 3394 2947 3432 2981
rect 3466 2947 3504 2981
rect 3538 2947 3576 2981
rect 3610 2947 3648 2981
rect 3682 2947 3720 2981
rect 3754 2947 3792 2981
rect 3826 2947 3864 2981
rect 3898 2947 3936 2981
rect 3970 2947 3983 2981
rect 68 2853 3983 2947
rect 68 2819 74 2853
rect 108 2819 386 2853
rect 420 2819 1084 2853
rect 1118 2819 1400 2853
rect 1434 2819 1616 2853
rect 1650 2819 1928 2853
rect 1962 2819 2240 2853
rect 2274 2819 2928 2853
rect 2962 2819 3983 2853
rect 68 2781 3983 2819
rect 68 2780 1400 2781
rect 68 2779 147 2780
tri 147 2779 148 2780 nw
tri 346 2779 347 2780 ne
rect 347 2779 459 2780
tri 459 2779 460 2780 nw
tri 1044 2779 1045 2780 ne
rect 1045 2779 1126 2780
rect 68 2776 116 2779
rect 68 2742 74 2776
rect 108 2748 116 2776
tri 116 2748 147 2779 nw
tri 347 2748 378 2779 ne
rect 378 2748 386 2779
rect 108 2742 114 2748
tri 114 2746 116 2748 nw
rect 68 2699 114 2742
rect 68 2665 74 2699
rect 108 2665 114 2699
rect 68 2622 114 2665
rect 68 2588 74 2622
rect 108 2588 114 2622
rect 68 2544 114 2588
rect 68 2510 74 2544
rect 108 2510 114 2544
rect 68 2466 114 2510
rect 68 2432 74 2466
rect 108 2432 114 2466
rect 68 2388 114 2432
rect 68 2354 74 2388
rect 108 2354 114 2388
rect 68 2310 114 2354
rect 68 2276 74 2310
rect 108 2276 114 2310
rect 68 2232 114 2276
rect 68 2198 74 2232
rect 108 2198 114 2232
rect 68 2154 114 2198
rect 68 2120 74 2154
rect 108 2120 114 2154
rect 68 2076 114 2120
rect 68 2042 74 2076
rect 108 2042 114 2076
rect 68 1998 114 2042
rect 68 1964 74 1998
rect 108 1964 114 1998
rect 68 1920 114 1964
rect 68 1886 74 1920
rect 108 1886 114 1920
rect 68 1874 114 1886
rect 224 2736 270 2748
tri 378 2746 380 2748 ne
rect 224 2702 230 2736
rect 264 2702 270 2736
rect 224 2661 270 2702
rect 224 2627 230 2661
rect 264 2627 270 2661
rect 224 2586 270 2627
rect 224 2552 230 2586
rect 264 2552 270 2586
rect 224 2511 270 2552
rect 224 2477 230 2511
rect 264 2477 270 2511
rect 224 2436 270 2477
rect 224 2402 230 2436
rect 264 2402 270 2436
rect 224 2361 270 2402
rect 224 2327 230 2361
rect 264 2327 270 2361
rect 224 2286 270 2327
rect 224 2252 230 2286
rect 264 2252 270 2286
rect 224 2211 270 2252
rect 224 2177 230 2211
rect 264 2177 270 2211
rect 224 2135 270 2177
rect 224 2101 230 2135
rect 264 2101 270 2135
rect 224 2059 270 2101
rect 224 2025 230 2059
rect 264 2025 270 2059
rect 224 1993 270 2025
rect 380 2745 386 2748
rect 420 2748 428 2779
tri 428 2748 459 2779 nw
tri 1045 2748 1076 2779 ne
rect 1076 2748 1084 2779
rect 420 2745 426 2748
tri 426 2746 428 2748 nw
rect 380 2705 426 2745
rect 380 2671 386 2705
rect 420 2671 426 2705
rect 380 2631 426 2671
rect 380 2597 386 2631
rect 420 2597 426 2631
rect 380 2557 426 2597
rect 380 2523 386 2557
rect 420 2523 426 2557
rect 380 2483 426 2523
rect 380 2449 386 2483
rect 420 2449 426 2483
rect 380 2409 426 2449
rect 380 2375 386 2409
rect 420 2375 426 2409
rect 380 2335 426 2375
rect 380 2301 386 2335
rect 420 2301 426 2335
rect 380 2261 426 2301
rect 380 2227 386 2261
rect 420 2227 426 2261
rect 380 2187 426 2227
rect 380 2153 386 2187
rect 420 2153 426 2187
rect 380 2113 426 2153
rect 380 2079 386 2113
rect 420 2079 426 2113
rect 380 2039 426 2079
rect 380 2005 386 2039
rect 420 2005 426 2039
tri 270 1993 272 1995 sw
rect 380 1993 426 2005
rect 490 2736 536 2748
rect 490 2702 496 2736
rect 530 2702 536 2736
rect 490 2661 536 2702
rect 490 2627 496 2661
rect 530 2627 536 2661
rect 490 2586 536 2627
rect 490 2552 496 2586
rect 530 2552 536 2586
rect 490 2511 536 2552
rect 490 2477 496 2511
rect 530 2477 536 2511
rect 490 2436 536 2477
rect 490 2402 496 2436
rect 530 2402 536 2436
rect 490 2361 536 2402
rect 490 2327 496 2361
rect 530 2327 536 2361
rect 490 2286 536 2327
rect 490 2252 496 2286
rect 530 2252 536 2286
rect 490 2211 536 2252
rect 490 2177 496 2211
rect 530 2177 536 2211
rect 490 2135 536 2177
rect 490 2101 496 2135
rect 530 2101 536 2135
rect 490 2059 536 2101
rect 490 2025 496 2059
rect 530 2025 536 2059
tri 488 1993 490 1995 se
rect 490 1993 536 2025
rect 224 1992 272 1993
tri 272 1992 273 1993 sw
tri 487 1992 488 1993 se
rect 488 1992 536 1993
rect 224 1983 273 1992
tri 273 1983 282 1992 sw
tri 478 1983 487 1992 se
rect 487 1983 536 1992
rect 224 1949 230 1983
rect 264 1961 282 1983
tri 282 1961 304 1983 sw
tri 456 1961 478 1983 se
rect 478 1961 496 1983
rect 264 1949 496 1961
rect 530 1949 536 1983
rect 224 1907 536 1949
rect 224 1873 230 1907
rect 264 1873 496 1907
rect 530 1873 536 1907
rect 224 1861 536 1873
rect 703 2736 755 2748
rect 703 2702 712 2736
rect 746 2702 755 2736
rect 703 2661 755 2702
rect 703 2627 712 2661
rect 746 2627 755 2661
rect 703 2586 755 2627
rect 703 2552 712 2586
rect 746 2552 755 2586
rect 703 2511 755 2552
rect 703 2477 712 2511
rect 746 2477 755 2511
rect 703 2436 755 2477
rect 703 2402 712 2436
rect 746 2402 755 2436
rect 703 2361 755 2402
rect 703 2327 712 2361
rect 746 2327 755 2361
rect 703 2286 755 2327
rect 703 2252 712 2286
rect 746 2252 755 2286
rect 703 2211 755 2252
rect 703 2177 712 2211
rect 746 2177 755 2211
rect 703 2173 755 2177
rect 703 2101 712 2121
rect 746 2101 755 2121
rect 703 2091 755 2101
rect 703 2025 712 2039
rect 746 2025 755 2039
rect 703 2008 755 2025
rect 703 1949 712 1956
rect 746 1949 755 1956
rect 703 1925 755 1949
rect 703 1861 755 1873
rect 922 2736 968 2748
tri 1076 2746 1078 2748 ne
rect 922 2702 928 2736
rect 962 2702 968 2736
rect 922 2661 968 2702
rect 922 2627 928 2661
rect 962 2627 968 2661
rect 922 2586 968 2627
rect 922 2552 928 2586
rect 962 2552 968 2586
rect 922 2511 968 2552
rect 922 2477 928 2511
rect 962 2477 968 2511
rect 922 2436 968 2477
rect 922 2402 928 2436
rect 962 2402 968 2436
rect 922 2361 968 2402
rect 922 2327 928 2361
rect 962 2327 968 2361
rect 922 2286 968 2327
rect 922 2252 928 2286
rect 962 2252 968 2286
rect 922 2211 968 2252
rect 922 2177 928 2211
rect 962 2177 968 2211
rect 922 2135 968 2177
rect 922 2101 928 2135
rect 962 2101 968 2135
rect 922 2059 968 2101
rect 922 2025 928 2059
rect 962 2025 968 2059
rect 922 1992 968 2025
rect 1078 2745 1084 2748
rect 1118 2748 1126 2779
tri 1126 2748 1158 2780 nw
tri 1360 2748 1392 2780 ne
rect 1392 2748 1400 2780
rect 1118 2747 1125 2748
tri 1125 2747 1126 2748 nw
rect 1118 2745 1124 2747
tri 1124 2746 1125 2747 nw
rect 1078 2705 1124 2745
rect 1078 2671 1084 2705
rect 1118 2671 1124 2705
rect 1078 2631 1124 2671
rect 1078 2597 1084 2631
rect 1118 2597 1124 2631
rect 1078 2557 1124 2597
rect 1078 2523 1084 2557
rect 1118 2523 1124 2557
rect 1078 2483 1124 2523
rect 1078 2449 1084 2483
rect 1118 2449 1124 2483
rect 1078 2409 1124 2449
rect 1078 2375 1084 2409
rect 1118 2375 1124 2409
rect 1078 2335 1124 2375
rect 1078 2301 1084 2335
rect 1118 2301 1124 2335
rect 1078 2261 1124 2301
rect 1078 2227 1084 2261
rect 1118 2227 1124 2261
rect 1078 2187 1124 2227
rect 1078 2153 1084 2187
rect 1118 2153 1124 2187
rect 1078 2112 1124 2153
rect 1078 2078 1084 2112
rect 1118 2078 1124 2112
rect 1078 2037 1124 2078
rect 1078 2003 1084 2037
rect 1118 2003 1124 2037
tri 968 1992 971 1995 sw
rect 922 1991 971 1992
tri 971 1991 972 1992 sw
rect 1078 1991 1124 2003
rect 1234 2736 1280 2748
tri 1392 2747 1393 2748 ne
rect 1393 2747 1400 2748
rect 1434 2780 1616 2781
rect 1434 2747 1441 2780
tri 1441 2747 1474 2780 nw
tri 1576 2747 1609 2780 ne
rect 1609 2747 1616 2780
rect 1650 2780 1928 2781
rect 1650 2748 1658 2780
tri 1658 2748 1690 2780 nw
tri 1888 2748 1920 2780 ne
rect 1920 2748 1928 2780
rect 1650 2747 1657 2748
tri 1657 2747 1658 2748 nw
tri 1393 2746 1394 2747 ne
rect 1234 2702 1240 2736
rect 1274 2702 1280 2736
rect 1234 2661 1280 2702
rect 1234 2627 1240 2661
rect 1274 2627 1280 2661
rect 1234 2586 1280 2627
rect 1234 2552 1240 2586
rect 1274 2552 1280 2586
rect 1234 2511 1280 2552
rect 1234 2477 1240 2511
rect 1274 2477 1280 2511
rect 1234 2436 1280 2477
rect 1234 2402 1240 2436
rect 1274 2402 1280 2436
rect 1234 2361 1280 2402
rect 1234 2327 1240 2361
rect 1274 2327 1280 2361
rect 1234 2286 1280 2327
rect 1234 2252 1240 2286
rect 1274 2252 1280 2286
rect 1234 2211 1280 2252
rect 1234 2177 1240 2211
rect 1274 2177 1280 2211
rect 1234 2135 1280 2177
rect 1234 2101 1240 2135
rect 1274 2101 1280 2135
rect 1234 2059 1280 2101
rect 1234 2025 1240 2059
rect 1274 2025 1280 2059
tri 1231 1992 1234 1995 se
rect 1234 1992 1280 2025
tri 1230 1991 1231 1992 se
rect 1231 1991 1280 1992
rect 922 1983 972 1991
tri 972 1983 980 1991 sw
tri 1222 1983 1230 1991 se
rect 1230 1983 1280 1991
rect 922 1949 928 1983
rect 962 1961 980 1983
tri 980 1961 1002 1983 sw
tri 1200 1961 1222 1983 se
rect 1222 1961 1240 1983
rect 962 1949 1240 1961
rect 1274 1949 1280 1983
rect 922 1907 1280 1949
rect 922 1873 928 1907
rect 962 1873 1240 1907
rect 1274 1873 1280 1907
rect 922 1861 1280 1873
rect 1394 2709 1440 2747
tri 1440 2746 1441 2747 nw
tri 1609 2746 1610 2747 ne
rect 1394 2675 1400 2709
rect 1434 2675 1440 2709
rect 1394 2637 1440 2675
rect 1394 2603 1400 2637
rect 1434 2603 1440 2637
rect 1394 2564 1440 2603
rect 1394 2530 1400 2564
rect 1434 2530 1440 2564
rect 1394 2491 1440 2530
rect 1394 2457 1400 2491
rect 1434 2457 1440 2491
rect 1394 2418 1440 2457
rect 1394 2384 1400 2418
rect 1434 2384 1440 2418
rect 1394 2345 1440 2384
rect 1394 2311 1400 2345
rect 1434 2311 1440 2345
rect 1394 2272 1440 2311
rect 1394 2238 1400 2272
rect 1434 2238 1440 2272
rect 1394 2199 1440 2238
rect 1394 2165 1400 2199
rect 1434 2165 1440 2199
rect 1394 2126 1440 2165
rect 1394 2092 1400 2126
rect 1434 2092 1440 2126
rect 1394 2053 1440 2092
rect 1394 2019 1400 2053
rect 1434 2019 1440 2053
rect 1394 1980 1440 2019
rect 1394 1946 1400 1980
rect 1434 1946 1440 1980
rect 1394 1907 1440 1946
rect 1394 1873 1400 1907
rect 1434 1873 1440 1907
rect 1394 1826 1440 1873
rect 1610 2709 1656 2747
tri 1656 2746 1657 2747 nw
rect 1610 2675 1616 2709
rect 1650 2675 1656 2709
rect 1610 2637 1656 2675
rect 1610 2603 1616 2637
rect 1650 2603 1656 2637
rect 1610 2564 1656 2603
rect 1610 2530 1616 2564
rect 1650 2530 1656 2564
rect 1610 2491 1656 2530
rect 1610 2457 1616 2491
rect 1650 2457 1656 2491
rect 1610 2418 1656 2457
rect 1610 2384 1616 2418
rect 1650 2384 1656 2418
rect 1610 2345 1656 2384
rect 1610 2311 1616 2345
rect 1650 2311 1656 2345
rect 1610 2272 1656 2311
rect 1610 2238 1616 2272
rect 1650 2238 1656 2272
rect 1610 2199 1656 2238
rect 1610 2165 1616 2199
rect 1650 2165 1656 2199
rect 1610 2126 1656 2165
rect 1610 2092 1616 2126
rect 1650 2092 1656 2126
rect 1610 2053 1656 2092
rect 1610 2019 1616 2053
rect 1650 2019 1656 2053
rect 1610 1980 1656 2019
rect 1610 1946 1616 1980
rect 1650 1946 1656 1980
rect 1610 1907 1656 1946
rect 1610 1873 1616 1907
rect 1650 1873 1656 1907
rect 1610 1861 1656 1873
rect 1763 2736 1815 2748
tri 1920 2747 1921 2748 ne
rect 1921 2747 1928 2748
rect 1962 2780 2240 2781
rect 1962 2748 1970 2780
tri 1970 2748 2002 2780 nw
tri 2200 2748 2232 2780 ne
rect 2232 2748 2240 2780
rect 1962 2747 1969 2748
tri 1969 2747 1970 2748 nw
tri 1921 2746 1922 2747 ne
rect 1763 2702 1772 2736
rect 1806 2702 1815 2736
rect 1763 2661 1815 2702
rect 1763 2627 1772 2661
rect 1806 2627 1815 2661
rect 1763 2586 1815 2627
rect 1763 2552 1772 2586
rect 1806 2552 1815 2586
rect 1763 2511 1815 2552
rect 1763 2477 1772 2511
rect 1806 2477 1815 2511
rect 1763 2436 1815 2477
rect 1763 2402 1772 2436
rect 1806 2402 1815 2436
rect 1763 2361 1815 2402
rect 1763 2327 1772 2361
rect 1806 2327 1815 2361
rect 1763 2286 1815 2327
rect 1763 2252 1772 2286
rect 1806 2252 1815 2286
rect 1763 2211 1815 2252
rect 1763 2177 1772 2211
rect 1806 2177 1815 2211
rect 1763 2166 1815 2177
rect 1763 2101 1772 2114
rect 1806 2101 1815 2114
rect 1763 2084 1815 2101
rect 1763 2025 1772 2032
rect 1806 2025 1815 2032
rect 1763 2002 1815 2025
rect 1763 1949 1772 1950
rect 1806 1949 1815 1950
rect 1763 1919 1815 1949
rect 1763 1861 1815 1867
rect 1922 2709 1968 2747
tri 1968 2746 1969 2747 nw
rect 1922 2675 1928 2709
rect 1962 2675 1968 2709
rect 1922 2637 1968 2675
rect 1922 2603 1928 2637
rect 1962 2603 1968 2637
rect 1922 2564 1968 2603
rect 1922 2530 1928 2564
rect 1962 2530 1968 2564
rect 1922 2491 1968 2530
rect 1922 2457 1928 2491
rect 1962 2457 1968 2491
rect 1922 2418 1968 2457
rect 1922 2384 1928 2418
rect 1962 2384 1968 2418
rect 1922 2345 1968 2384
rect 1922 2311 1928 2345
rect 1962 2311 1968 2345
rect 1922 2272 1968 2311
rect 1922 2238 1928 2272
rect 1962 2238 1968 2272
rect 1922 2199 1968 2238
rect 1922 2165 1928 2199
rect 1962 2165 1968 2199
rect 1922 2126 1968 2165
rect 1922 2092 1928 2126
rect 1962 2092 1968 2126
rect 1922 2053 1968 2092
rect 1922 2019 1928 2053
rect 1962 2019 1968 2053
rect 1922 1980 1968 2019
rect 1922 1946 1928 1980
rect 1962 1946 1968 1980
rect 1922 1907 1968 1946
rect 1922 1873 1928 1907
rect 1962 1873 1968 1907
rect 1922 1861 1968 1873
rect 2075 2736 2127 2748
tri 2232 2747 2233 2748 ne
rect 2233 2747 2240 2748
rect 2274 2780 3983 2781
rect 2274 2776 2310 2780
tri 2310 2776 2314 2780 nw
tri 2888 2776 2892 2780 ne
rect 2892 2776 2970 2780
rect 2274 2748 2282 2776
tri 2282 2748 2310 2776 nw
tri 2892 2748 2920 2776 ne
rect 2920 2748 2928 2776
rect 2274 2747 2280 2748
tri 2233 2746 2234 2747 ne
rect 2075 2702 2084 2736
rect 2118 2702 2127 2736
rect 2075 2661 2127 2702
rect 2075 2627 2084 2661
rect 2118 2627 2127 2661
rect 2075 2586 2127 2627
rect 2075 2552 2084 2586
rect 2118 2552 2127 2586
rect 2075 2511 2127 2552
rect 2075 2477 2084 2511
rect 2118 2477 2127 2511
rect 2075 2436 2127 2477
rect 2075 2402 2084 2436
rect 2118 2402 2127 2436
rect 2075 2361 2127 2402
rect 2075 2327 2084 2361
rect 2118 2327 2127 2361
rect 2075 2286 2127 2327
rect 2075 2252 2084 2286
rect 2118 2252 2127 2286
rect 2075 2211 2127 2252
rect 2075 2177 2084 2211
rect 2118 2177 2127 2211
rect 2075 2166 2127 2177
rect 2075 2101 2084 2114
rect 2118 2101 2127 2114
rect 2075 2084 2127 2101
rect 2075 2025 2084 2032
rect 2118 2025 2127 2032
rect 2075 2002 2127 2025
rect 2075 1949 2084 1950
rect 2118 1949 2127 1950
rect 2075 1919 2127 1949
rect 2075 1861 2127 1867
rect 2234 2709 2280 2747
tri 2280 2746 2282 2748 nw
rect 2234 2675 2240 2709
rect 2274 2675 2280 2709
rect 2234 2637 2280 2675
rect 2234 2603 2240 2637
rect 2274 2603 2280 2637
rect 2234 2564 2280 2603
rect 2234 2530 2240 2564
rect 2274 2530 2280 2564
rect 2234 2491 2280 2530
rect 2234 2457 2240 2491
rect 2274 2457 2280 2491
rect 2234 2418 2280 2457
rect 2234 2384 2240 2418
rect 2274 2384 2280 2418
rect 2234 2345 2280 2384
rect 2234 2311 2240 2345
rect 2274 2311 2280 2345
rect 2234 2272 2280 2311
rect 2234 2238 2240 2272
rect 2274 2238 2280 2272
rect 2234 2199 2280 2238
rect 2234 2165 2240 2199
rect 2274 2165 2280 2199
rect 2234 2126 2280 2165
rect 2234 2092 2240 2126
rect 2274 2092 2280 2126
rect 2234 2053 2280 2092
rect 2234 2019 2240 2053
rect 2274 2019 2280 2053
rect 2234 1980 2280 2019
rect 2234 1946 2240 1980
rect 2274 1946 2280 1980
rect 2234 1907 2280 1946
rect 2234 1873 2240 1907
rect 2274 1873 2280 1907
rect 2234 1861 2280 1873
rect 2390 2736 2436 2748
rect 2390 2702 2396 2736
rect 2430 2702 2436 2736
rect 2390 2661 2436 2702
rect 2390 2627 2396 2661
rect 2430 2627 2436 2661
rect 2390 2586 2436 2627
rect 2390 2552 2396 2586
rect 2430 2552 2436 2586
rect 2390 2511 2436 2552
rect 2390 2477 2396 2511
rect 2430 2477 2436 2511
rect 2390 2436 2436 2477
rect 2390 2402 2396 2436
rect 2430 2402 2436 2436
rect 2766 2736 2812 2748
tri 2920 2746 2922 2748 ne
rect 2766 2702 2772 2736
rect 2806 2702 2812 2736
rect 2766 2658 2812 2702
rect 2766 2624 2772 2658
rect 2806 2624 2812 2658
rect 2766 2580 2812 2624
rect 2766 2546 2772 2580
rect 2806 2546 2812 2580
rect 2766 2502 2812 2546
rect 2766 2468 2772 2502
rect 2806 2468 2812 2502
rect 2766 2424 2812 2468
rect 2390 2390 2436 2402
tri 2436 2390 2458 2412 sw
rect 2766 2390 2772 2424
rect 2806 2390 2812 2424
rect 2390 2387 2458 2390
tri 2458 2387 2461 2390 sw
rect 2390 2378 2461 2387
tri 2461 2378 2470 2387 sw
rect 2390 2366 2546 2378
rect 2390 2361 2506 2366
rect 2390 2327 2396 2361
rect 2430 2332 2506 2361
rect 2540 2332 2546 2366
rect 2430 2327 2546 2332
rect 2390 2286 2546 2327
rect 2390 2252 2396 2286
rect 2430 2281 2546 2286
rect 2430 2252 2506 2281
rect 2390 2247 2506 2252
rect 2540 2247 2546 2281
rect 2390 2211 2546 2247
rect 2390 2177 2396 2211
rect 2430 2196 2546 2211
rect 2430 2177 2506 2196
rect 2390 2162 2506 2177
rect 2540 2162 2546 2196
rect 2390 2135 2546 2162
rect 2390 2101 2396 2135
rect 2430 2111 2546 2135
rect 2430 2101 2506 2111
rect 2390 2077 2506 2101
rect 2540 2077 2546 2111
rect 2390 2059 2546 2077
rect 2390 2025 2396 2059
rect 2430 2026 2546 2059
rect 2430 2025 2506 2026
rect 2390 1992 2506 2025
rect 2540 1992 2546 2026
rect 2390 1983 2546 1992
rect 2390 1949 2396 1983
rect 2430 1949 2546 1983
rect 2390 1941 2546 1949
rect 2390 1907 2506 1941
rect 2540 1907 2546 1941
rect 2390 1873 2396 1907
rect 2430 1895 2546 1907
rect 2656 2366 2702 2378
rect 2656 2332 2662 2366
rect 2696 2332 2702 2366
rect 2656 2281 2702 2332
rect 2656 2247 2662 2281
rect 2696 2247 2702 2281
rect 2656 2196 2702 2247
rect 2656 2162 2662 2196
rect 2696 2162 2702 2196
rect 2656 2111 2702 2162
rect 2656 2077 2662 2111
rect 2696 2077 2702 2111
rect 2656 2026 2702 2077
rect 2656 1992 2662 2026
rect 2696 1992 2702 2026
rect 2656 1941 2702 1992
rect 2656 1907 2662 1941
rect 2696 1907 2702 1941
rect 2430 1873 2436 1895
rect 2390 1861 2436 1873
tri 2436 1861 2470 1895 nw
tri 1440 1826 1471 1857 sw
rect 2656 1826 2702 1907
rect 2766 2346 2812 2390
rect 2766 2312 2772 2346
rect 2806 2312 2812 2346
rect 2766 2267 2812 2312
rect 2766 2233 2772 2267
rect 2806 2233 2812 2267
rect 2766 2188 2812 2233
rect 2766 2154 2772 2188
rect 2806 2154 2812 2188
rect 2766 2109 2812 2154
rect 2766 2075 2772 2109
rect 2806 2075 2812 2109
rect 2766 2030 2812 2075
rect 2766 1996 2772 2030
rect 2806 1996 2812 2030
rect 2766 1909 2812 1996
rect 2922 2742 2928 2748
rect 2962 2748 2970 2776
tri 2970 2748 3002 2780 nw
rect 2962 2742 2968 2748
tri 2968 2746 2970 2748 nw
rect 2922 2699 2968 2742
rect 2922 2665 2928 2699
rect 2962 2665 2968 2699
rect 2922 2621 2968 2665
rect 2922 2587 2928 2621
rect 2962 2587 2968 2621
rect 2922 2543 2968 2587
rect 2922 2509 2928 2543
rect 2962 2509 2968 2543
rect 2922 2465 2968 2509
rect 2922 2431 2928 2465
rect 2962 2431 2968 2465
rect 2922 2387 2968 2431
rect 2922 2353 2928 2387
rect 2962 2353 2968 2387
rect 2922 2309 2968 2353
rect 2922 2275 2928 2309
rect 2962 2275 2968 2309
rect 2922 2231 2968 2275
rect 2922 2197 2928 2231
rect 2962 2197 2968 2231
rect 2922 2153 2968 2197
rect 2922 2119 2928 2153
rect 2962 2119 2968 2153
rect 2922 2075 2968 2119
rect 2922 2041 2928 2075
rect 2962 2041 2968 2075
rect 2922 1997 2968 2041
rect 2922 1963 2928 1997
rect 2962 1963 2968 1997
rect 2922 1951 2968 1963
rect 3078 2736 3124 2748
rect 3078 2702 3084 2736
rect 3118 2702 3124 2736
rect 3078 2661 3124 2702
rect 3078 2627 3084 2661
rect 3118 2627 3124 2661
rect 3078 2586 3124 2627
rect 3078 2552 3084 2586
rect 3118 2552 3124 2586
rect 3078 2511 3124 2552
rect 3078 2477 3084 2511
rect 3118 2477 3124 2511
rect 3078 2436 3124 2477
rect 3078 2402 3084 2436
rect 3118 2402 3124 2436
rect 3078 2361 3124 2402
rect 3446 2439 3831 2445
rect 3446 2405 3458 2439
rect 3492 2405 3530 2439
rect 3564 2405 3831 2439
rect 3446 2399 3831 2405
tri 3751 2371 3779 2399 ne
rect 3779 2371 3831 2399
rect 3078 2327 3084 2361
rect 3118 2327 3124 2361
rect 3078 2286 3124 2327
rect 3637 2365 3689 2371
tri 3779 2365 3785 2371 ne
rect 3078 2252 3084 2286
rect 3118 2252 3124 2286
rect 3384 2253 3392 2305
rect 3444 2253 3456 2305
rect 3508 2253 3514 2305
rect 3637 2301 3689 2313
rect 3785 2337 3791 2371
rect 3825 2337 3831 2371
rect 3785 2299 3831 2337
rect 3785 2265 3791 2299
rect 3825 2265 3831 2299
rect 3785 2253 3831 2265
rect 3885 2364 3937 2370
rect 3885 2300 3937 2312
rect 3078 2211 3124 2252
rect 3637 2241 3689 2249
rect 3885 2240 3937 2248
rect 3078 2177 3084 2211
rect 3118 2177 3124 2211
rect 3078 2136 3124 2177
rect 3078 2102 3084 2136
rect 3118 2102 3124 2136
rect 3078 2060 3124 2102
rect 3078 2026 3084 2060
rect 3118 2026 3124 2060
rect 3078 1984 3124 2026
rect 3078 1950 3084 1984
rect 3118 1950 3124 1984
tri 2812 1909 2846 1943 sw
rect 3078 1938 3124 1950
rect 3601 2154 3721 2160
rect 3653 2102 3669 2154
rect 3601 2079 3721 2102
rect 3653 2027 3669 2079
rect 3601 2003 3721 2027
rect 3653 1951 3669 2003
tri 3124 1938 3134 1948 sw
rect 3601 1945 3721 1951
rect 3078 1928 3134 1938
tri 3134 1928 3144 1938 sw
tri 3078 1909 3097 1928 ne
rect 3097 1909 3144 1928
rect 2766 1904 2980 1909
tri 2980 1904 2985 1909 sw
tri 3097 1904 3102 1909 ne
rect 3102 1904 3144 1909
rect 2766 1868 2985 1904
tri 2985 1868 3021 1904 sw
rect 2766 1863 3021 1868
tri 2941 1860 2944 1863 ne
rect 2944 1860 3021 1863
tri 3102 1862 3144 1904 ne
tri 3144 1862 3210 1928 sw
tri 3144 1860 3146 1862 ne
rect 3146 1860 3210 1862
tri 2702 1826 2736 1860 sw
tri 2944 1829 2975 1860 ne
rect 2975 1826 3021 1860
tri 3021 1826 3055 1860 sw
tri 3146 1826 3180 1860 ne
rect 3180 1842 3210 1860
tri 3210 1842 3230 1862 sw
rect 3180 1826 3236 1842
rect 125 1773 131 1825
rect 183 1773 195 1825
rect 247 1817 370 1825
rect 265 1783 324 1817
rect 358 1783 370 1817
rect 247 1773 370 1783
rect 543 1774 549 1826
rect 601 1817 613 1826
rect 665 1817 902 1826
rect 612 1783 613 1817
rect 684 1783 784 1817
rect 818 1783 856 1817
rect 890 1783 902 1817
rect 601 1774 613 1783
rect 665 1774 902 1783
rect 973 1817 1042 1826
rect 1094 1817 1106 1826
rect 1158 1817 1229 1826
rect 973 1783 985 1817
rect 1019 1783 1042 1817
rect 1158 1783 1183 1817
rect 1217 1783 1229 1817
rect 973 1774 1042 1783
rect 1094 1774 1106 1783
rect 1158 1774 1229 1783
rect 1394 1825 1471 1826
tri 1471 1825 1472 1826 sw
rect 1394 1823 1472 1825
tri 1472 1823 1474 1825 sw
rect 1394 1817 1525 1823
rect 1394 1783 1407 1817
rect 1441 1783 1479 1817
rect 1513 1783 1525 1817
rect 1394 1777 1525 1783
rect 1557 1773 1563 1825
rect 1615 1773 1627 1825
rect 1679 1817 1906 1825
rect 1707 1783 1767 1817
rect 1801 1783 1860 1817
rect 1894 1783 1906 1817
rect 1679 1773 1906 1783
rect 1980 1817 2290 1825
rect 1980 1783 1992 1817
rect 2026 1783 2086 1817
rect 2120 1783 2179 1817
rect 2213 1783 2290 1817
rect 1980 1773 2290 1783
rect 2342 1773 2354 1825
rect 2406 1817 2424 1825
rect 2412 1783 2424 1817
rect 2406 1773 2424 1783
rect 2498 1774 2506 1826
rect 2558 1774 2570 1826
rect 2622 1774 2628 1826
rect 2656 1774 2791 1826
rect 2843 1774 2855 1826
rect 2907 1774 2913 1826
rect 2975 1774 2981 1826
rect 3033 1774 3045 1826
rect 3097 1774 3105 1826
tri 3180 1823 3183 1826 ne
rect 3183 1823 3236 1826
tri 3183 1796 3210 1823 ne
rect 3210 1796 3236 1823
tri 3210 1790 3216 1796 ne
rect 3216 1790 3236 1796
rect 3288 1790 3300 1842
rect 3352 1790 3358 1842
rect 91 1673 131 1725
rect 183 1673 195 1725
rect 247 1673 2290 1725
rect 2342 1673 2354 1725
rect 2406 1673 3392 1725
rect 3444 1673 3456 1725
rect 3508 1673 4883 1725
rect 4935 1673 4947 1725
rect 4999 1673 5503 1725
rect 1036 1513 1042 1565
rect 1094 1513 1106 1565
rect 1158 1513 1563 1565
rect 1615 1513 1627 1565
rect 1679 1513 3891 1565
rect 3943 1513 3955 1565
rect 4007 1513 4013 1565
rect 254 1433 1192 1485
rect 1244 1433 1256 1485
rect 1308 1433 4293 1485
rect 4345 1433 4357 1485
rect 4409 1433 4415 1485
rect 703 1353 709 1405
rect 761 1353 773 1405
rect 825 1353 2506 1405
rect 2558 1353 2570 1405
rect 2622 1353 2728 1405
rect 2780 1353 2792 1405
rect 2844 1353 4576 1405
rect 4628 1353 4640 1405
rect 4692 1353 4774 1405
rect 1713 1273 1719 1325
rect 1771 1273 1783 1325
rect 1835 1273 2594 1325
rect 2646 1273 2658 1325
rect 2710 1273 2716 1325
rect 2075 1193 2081 1245
rect 2133 1193 2145 1245
rect 2197 1193 4470 1245
rect 4522 1193 4534 1245
rect 4586 1193 4592 1245
rect 254 1109 3767 1161
rect 3819 1109 3831 1161
rect 3883 1109 3889 1161
rect 3230 796 3236 848
rect 3288 796 3300 848
rect 3352 796 5636 848
rect 5688 796 5700 848
rect 5752 796 5758 848
rect 2975 678 2981 730
rect 3033 678 3045 730
rect 3097 678 5480 730
rect 5532 678 5544 730
rect 5596 678 5602 730
rect 2878 644 5377 650
rect 2930 598 5377 644
rect 5429 598 5441 650
rect 5493 598 5499 650
rect 2878 580 2930 592
tri 2930 564 2964 598 nw
rect 2878 522 2930 528
rect 4459 547 4511 553
tri 4425 477 4459 511 se
rect 4459 483 4511 495
rect 254 431 4459 477
rect 254 425 4511 431
rect 254 333 549 385
rect 601 333 613 385
rect 665 333 1875 385
rect 1927 333 1939 385
rect 1991 333 3652 385
tri 3427 299 3461 333 ne
rect 100 280 549 289
rect 601 280 613 289
rect 665 280 1080 289
rect 100 246 112 280
rect 146 246 189 280
rect 223 246 266 280
rect 300 246 343 280
rect 377 246 420 280
rect 454 246 497 280
rect 531 246 549 280
rect 608 246 613 280
rect 685 246 728 280
rect 762 246 805 280
rect 839 246 882 280
rect 916 246 958 280
rect 992 246 1034 280
rect 1068 246 1080 280
rect 100 237 549 246
rect 601 237 613 246
rect 665 237 1080 246
rect 1186 237 1192 289
rect 1244 237 1258 289
rect 1310 237 1316 289
rect 1403 280 1875 289
rect 1403 246 1415 280
rect 1449 246 1492 280
rect 1526 246 1569 280
rect 1603 246 1646 280
rect 1680 246 1723 280
rect 1757 246 1800 280
rect 1834 246 1875 280
rect 1403 237 1875 246
rect 1927 237 1939 289
rect 1991 280 2383 289
rect 1991 246 2031 280
rect 2065 246 2108 280
rect 2142 246 2185 280
rect 2219 246 2261 280
rect 2295 246 2337 280
rect 2371 246 2383 280
rect 1991 237 2383 246
rect 2495 280 2804 289
rect 2495 246 2507 280
rect 2541 246 2585 280
rect 2619 246 2663 280
rect 2697 246 2741 280
rect 2775 246 2804 280
rect 2495 237 2804 246
rect 2856 237 2868 289
rect 2920 280 3250 289
rect 2930 246 2973 280
rect 3007 246 3050 280
rect 3084 246 3127 280
rect 3161 246 3204 280
rect 3238 246 3250 280
rect 2920 237 3250 246
rect 3461 280 3591 333
tri 3591 299 3625 333 nw
rect 4477 289 5195 291
rect 3461 246 3473 280
rect 3507 246 3545 280
rect 3579 246 3591 280
rect 3461 240 3591 246
rect 3787 237 3795 289
rect 3847 237 3859 289
rect 3911 237 3917 289
rect 4113 280 4183 289
rect 4113 246 4125 280
rect 4159 246 4183 280
rect 4113 237 4183 246
rect 4235 237 4247 289
rect 4299 237 4305 289
rect 4477 285 4652 289
rect 4704 285 4716 289
rect 4768 285 5195 289
rect 4477 251 4489 285
rect 4523 251 4562 285
rect 4596 251 4635 285
rect 4704 251 4708 285
rect 4768 251 4781 285
rect 4815 251 4854 285
rect 4888 251 4926 285
rect 4960 251 4998 285
rect 5032 251 5070 285
rect 5104 251 5142 285
rect 5176 251 5195 285
rect 4477 239 4652 251
tri 4644 237 4646 239 ne
rect 4646 237 4652 239
rect 4704 237 4716 251
rect 4768 239 5195 251
rect 5247 239 5259 291
rect 5311 239 5317 291
rect 5348 280 5377 292
rect 5429 280 5441 292
rect 5348 246 5360 280
rect 5429 246 5433 280
rect 5348 240 5377 246
rect 5429 240 5441 246
rect 5493 240 5499 292
rect 4768 237 4774 239
tri 4774 237 4776 239 nw
rect 5550 237 5556 289
rect 5608 280 5620 289
rect 5672 280 5695 289
rect 5611 246 5620 280
rect 5683 246 5695 280
rect 5608 237 5620 246
rect 5672 237 5695 246
tri 5541 208 5550 217 se
rect 5550 208 5611 237
rect 38 196 84 208
rect 38 162 44 196
rect 78 162 84 196
rect 38 122 84 162
rect 38 88 44 122
rect 78 88 84 122
rect 38 48 84 88
rect 38 14 44 48
rect 78 14 84 48
rect 38 -26 84 14
rect 38 -60 44 -26
rect 78 -60 84 -26
rect 38 -100 84 -60
rect 38 -134 44 -100
rect 78 -134 84 -100
rect 38 -174 84 -134
rect 38 -208 44 -174
rect 78 -208 84 -174
rect 38 -248 84 -208
rect 38 -282 44 -248
rect 78 -282 84 -248
rect 38 -322 84 -282
rect 38 -356 44 -322
rect 78 -356 84 -322
rect 38 -395 84 -356
rect 38 -429 44 -395
rect 78 -429 84 -395
rect 38 -468 84 -429
rect 38 -502 44 -468
rect 78 -502 84 -468
rect 38 -541 84 -502
rect 38 -575 44 -541
rect 78 -575 84 -541
rect -467 -638 -461 -586
rect -409 -638 -376 -586
rect -324 -638 -291 -586
rect -239 -638 -207 -586
rect -155 -638 -123 -586
rect -71 -638 -65 -586
rect -467 -696 -65 -638
rect -467 -748 -461 -696
rect -409 -748 -376 -696
rect -324 -748 -291 -696
rect -239 -748 -207 -696
rect -155 -748 -123 -696
rect -71 -748 -65 -696
rect 38 -614 84 -575
rect 38 -648 44 -614
rect 78 -648 84 -614
rect 38 -674 84 -648
rect 254 196 5276 208
rect 254 162 260 196
rect 294 162 692 196
rect 726 162 1124 196
rect 1158 162 1556 196
rect 1590 162 1988 196
rect 2022 162 2420 196
rect 2454 162 2852 196
rect 2886 162 3284 196
rect 3318 162 3394 196
rect 3428 162 4372 196
rect 4406 162 4804 196
rect 4838 162 5236 196
rect 5270 162 5276 196
tri 5516 183 5541 208 se
rect 5541 183 5611 208
tri 5611 203 5645 237 nw
rect 254 124 5276 162
tri 5373 137 5419 183 se
rect 5419 137 5611 183
rect 254 121 4372 124
rect 254 87 260 121
rect 294 108 692 121
rect 294 87 395 108
tri 395 87 416 108 nw
tri 623 87 644 108 ne
rect 644 87 692 108
rect 726 108 1124 121
rect 726 87 777 108
tri 777 87 798 108 nw
tri 1055 103 1060 108 ne
rect 1060 103 1124 108
tri 1060 87 1076 103 ne
rect 1076 87 1124 103
rect 1158 108 1556 121
rect 1158 106 1228 108
tri 1228 106 1230 108 nw
tri 1487 106 1489 108 ne
rect 1489 106 1556 108
rect 1158 87 1209 106
tri 1209 87 1228 106 nw
tri 1489 103 1492 106 ne
rect 1492 103 1556 106
tri 1492 87 1508 103 ne
rect 1508 87 1556 103
rect 1590 108 1988 121
rect 1590 106 1660 108
tri 1660 106 1662 108 nw
tri 1919 106 1921 108 ne
rect 1921 106 1988 108
rect 1590 87 1641 106
tri 1641 87 1660 106 nw
tri 1921 103 1924 106 ne
rect 1924 103 1988 106
tri 1924 87 1940 103 ne
rect 1940 87 1988 103
rect 2022 108 2420 121
rect 2022 106 2092 108
tri 2092 106 2094 108 nw
tri 2351 106 2353 108 ne
rect 2353 106 2420 108
rect 2022 87 2073 106
tri 2073 87 2092 106 nw
tri 2353 103 2356 106 ne
rect 2356 103 2420 106
tri 2356 87 2372 103 ne
rect 2372 87 2420 103
rect 2454 108 2852 121
rect 2454 106 2524 108
tri 2524 106 2526 108 nw
tri 2783 106 2785 108 ne
rect 2785 106 2852 108
rect 2454 87 2505 106
tri 2505 87 2524 106 nw
tri 2785 103 2788 106 ne
rect 2788 103 2852 106
tri 2788 87 2804 103 ne
rect 2804 87 2852 103
rect 2886 108 3284 121
rect 2886 106 2956 108
tri 2956 106 2958 108 nw
tri 3244 106 3246 108 ne
rect 3246 106 3284 108
rect 2886 87 2937 106
tri 2937 87 2956 106 nw
tri 3246 87 3265 106 ne
rect 3265 87 3284 106
rect 3318 87 3394 121
rect 3428 108 4372 121
rect 3428 90 3450 108
tri 3450 90 3468 108 nw
tri 4336 90 4354 108 ne
rect 4354 90 4372 108
rect 4406 108 4804 124
rect 4406 90 4424 108
tri 4424 90 4442 108 nw
tri 4768 90 4786 108 ne
rect 4786 90 4804 108
rect 4838 108 5236 124
rect 4838 90 4856 108
tri 4856 90 4874 108 nw
tri 5200 90 5218 108 ne
rect 5218 90 5236 108
rect 5270 90 5276 124
rect 3428 87 3438 90
rect 254 79 387 87
tri 387 79 395 87 nw
tri 644 79 652 87 ne
rect 652 79 766 87
rect 254 76 384 79
tri 384 76 387 79 nw
tri 652 76 655 79 ne
rect 655 76 766 79
tri 766 76 777 87 nw
tri 1076 76 1087 87 ne
rect 1087 76 1198 87
tri 1198 76 1209 87 nw
tri 1508 76 1519 87 ne
rect 1519 76 1630 87
tri 1630 76 1641 87 nw
tri 1940 76 1951 87 ne
rect 1951 76 2062 87
tri 2062 76 2073 87 nw
tri 2372 76 2383 87 ne
rect 2383 76 2494 87
tri 2494 76 2505 87 nw
tri 2804 76 2815 87 ne
rect 2815 76 2926 87
tri 2926 76 2937 87 nw
tri 3265 76 3276 87 ne
rect 3276 78 3438 87
tri 3438 78 3450 90 nw
tri 4354 78 4366 90 ne
rect 4366 78 4412 90
tri 4412 78 4424 90 nw
tri 4786 78 4798 90 ne
rect 4798 78 4844 90
tri 4844 78 4856 90 nw
tri 5218 78 5230 90 ne
rect 5230 78 5276 90
tri 5356 120 5373 137 se
rect 5373 120 5411 137
rect 5356 109 5411 120
tri 5411 109 5439 137 nw
rect 5666 109 5718 121
rect 5356 108 5410 109
tri 5410 108 5411 109 nw
rect 3276 76 3436 78
tri 3436 76 3438 78 nw
rect 254 75 383 76
tri 383 75 384 76 nw
rect 254 46 373 75
tri 373 65 383 75 nw
rect 254 12 260 46
rect 294 12 373 46
rect 254 -29 373 12
rect 254 -63 260 -29
rect 294 -63 373 -29
rect 254 -104 373 -63
rect 254 -138 260 -104
rect 294 -138 373 -104
rect 254 -179 373 -138
rect 254 -213 260 -179
rect 294 -213 373 -179
rect 254 -254 373 -213
rect 254 -288 260 -254
rect 294 -288 373 -254
rect 254 -329 373 -288
rect 254 -363 260 -329
rect 294 -363 373 -329
rect 254 -404 373 -363
rect 254 -438 260 -404
rect 294 -438 373 -404
rect 254 -479 373 -438
rect 254 -513 260 -479
rect 294 -513 373 -479
rect 254 -554 373 -513
rect 254 -588 260 -554
rect 294 -588 373 -554
rect 254 -628 373 -588
rect 254 -662 260 -628
rect 294 -662 373 -628
tri 84 -674 86 -672 sw
rect 254 -674 373 -662
rect 444 64 551 76
tri 655 75 656 76 ne
rect 656 75 765 76
tri 765 75 766 76 nw
tri 656 74 657 75 ne
rect 444 30 476 64
rect 510 30 551 64
rect 444 -11 551 30
rect 444 -45 476 -11
rect 510 -45 551 -11
rect 444 -86 551 -45
rect 444 -120 476 -86
rect 510 -120 551 -86
rect 444 -161 551 -120
rect 444 -195 476 -161
rect 510 -195 551 -161
rect 444 -236 551 -195
rect 444 -270 476 -236
rect 510 -270 551 -236
rect 444 -311 551 -270
rect 444 -345 476 -311
rect 510 -345 551 -311
rect 444 -386 551 -345
rect 444 -420 476 -386
rect 510 -420 551 -386
rect 444 -461 551 -420
rect 444 -495 476 -461
rect 510 -495 551 -461
rect 444 -536 551 -495
rect 444 -570 476 -536
rect 510 -570 551 -536
rect 444 -611 551 -570
rect 444 -645 476 -611
rect 510 -645 551 -611
tri 442 -674 444 -672 se
rect 444 -674 551 -645
rect 657 46 764 75
tri 764 74 765 75 nw
rect 657 12 692 46
rect 726 12 764 46
rect 657 -29 764 12
rect 657 -63 692 -29
rect 726 -63 764 -29
rect 657 -104 764 -63
rect 657 -138 692 -104
rect 726 -138 764 -104
rect 657 -179 764 -138
rect 657 -213 692 -179
rect 726 -213 764 -179
rect 657 -254 764 -213
rect 657 -288 692 -254
rect 726 -288 764 -254
rect 657 -329 764 -288
rect 657 -363 692 -329
rect 726 -363 764 -329
rect 657 -404 764 -363
rect 657 -438 692 -404
rect 726 -438 764 -404
rect 657 -479 764 -438
rect 657 -513 692 -479
rect 726 -513 764 -479
rect 657 -554 764 -513
rect 657 -588 692 -554
rect 726 -588 764 -554
rect 657 -628 764 -588
rect 657 -662 692 -628
rect 726 -662 764 -628
rect 827 70 956 76
tri 1087 75 1088 76 ne
rect 1088 75 1197 76
tri 1197 75 1198 76 nw
tri 1088 74 1089 75 ne
rect 879 18 903 70
rect 955 18 956 70
rect 827 -11 956 18
rect 827 -19 908 -11
rect 942 -19 956 -11
rect 879 -71 903 -19
rect 955 -71 956 -19
rect 827 -86 956 -71
rect 827 -108 908 -86
rect 942 -108 956 -86
rect 879 -160 903 -108
rect 955 -160 956 -108
rect 827 -161 956 -160
rect 827 -195 908 -161
rect 942 -195 956 -161
rect 827 -197 956 -195
rect 879 -249 903 -197
rect 955 -249 956 -197
rect 827 -270 908 -249
rect 942 -270 956 -249
rect 827 -311 956 -270
rect 827 -345 908 -311
rect 942 -345 956 -311
rect 827 -386 956 -345
rect 827 -420 908 -386
rect 942 -420 956 -386
rect 827 -461 956 -420
rect 827 -495 908 -461
rect 942 -495 956 -461
rect 827 -536 956 -495
rect 827 -570 908 -536
rect 942 -570 956 -536
rect 827 -611 956 -570
rect 827 -645 908 -611
rect 942 -645 956 -611
tri 821 -662 827 -656 se
rect 827 -662 956 -645
tri 551 -674 553 -672 sw
rect 657 -674 764 -662
tri 809 -674 821 -662 se
rect 821 -674 956 -662
rect 1089 46 1196 75
tri 1196 74 1197 75 nw
rect 1089 12 1124 46
rect 1158 12 1196 46
rect 1089 -29 1196 12
rect 1089 -63 1124 -29
rect 1158 -63 1196 -29
rect 1089 -104 1196 -63
rect 1089 -138 1124 -104
rect 1158 -138 1196 -104
rect 1089 -179 1196 -138
rect 1089 -213 1124 -179
rect 1158 -213 1196 -179
rect 1089 -254 1196 -213
rect 1089 -288 1124 -254
rect 1158 -288 1196 -254
rect 1089 -329 1196 -288
rect 1089 -363 1124 -329
rect 1158 -363 1196 -329
rect 1089 -404 1196 -363
rect 1089 -438 1124 -404
rect 1158 -438 1196 -404
rect 1089 -479 1196 -438
rect 1089 -513 1124 -479
rect 1158 -513 1196 -479
rect 1089 -554 1196 -513
rect 1089 -588 1124 -554
rect 1158 -588 1196 -554
rect 1089 -628 1196 -588
rect 1089 -662 1124 -628
rect 1158 -662 1196 -628
rect 1089 -674 1196 -662
rect 1308 64 1415 76
tri 1519 75 1520 76 ne
rect 1520 75 1629 76
tri 1629 75 1630 76 nw
tri 1520 74 1521 75 ne
rect 1308 30 1340 64
rect 1374 30 1415 64
rect 1308 -11 1415 30
rect 1308 -45 1340 -11
rect 1374 -45 1415 -11
rect 1308 -86 1415 -45
rect 1308 -120 1340 -86
rect 1374 -120 1415 -86
rect 1308 -161 1415 -120
rect 1308 -195 1340 -161
rect 1374 -195 1415 -161
rect 1308 -236 1415 -195
rect 1308 -270 1340 -236
rect 1374 -270 1415 -236
rect 1308 -311 1415 -270
rect 1308 -345 1340 -311
rect 1374 -345 1415 -311
rect 1308 -386 1415 -345
rect 1308 -420 1340 -386
rect 1374 -420 1415 -386
rect 1308 -461 1415 -420
rect 1308 -495 1340 -461
rect 1374 -495 1415 -461
rect 1308 -536 1415 -495
rect 1308 -570 1340 -536
rect 1374 -570 1415 -536
rect 1308 -611 1415 -570
rect 1308 -645 1340 -611
rect 1374 -645 1415 -611
rect 1308 -674 1415 -645
rect 1521 46 1628 75
tri 1628 74 1629 75 nw
rect 1521 12 1556 46
rect 1590 12 1628 46
rect 1521 -29 1628 12
rect 1521 -63 1556 -29
rect 1590 -63 1628 -29
rect 1521 -104 1628 -63
rect 1521 -138 1556 -104
rect 1590 -138 1628 -104
rect 1521 -179 1628 -138
rect 1521 -213 1556 -179
rect 1590 -213 1628 -179
rect 1521 -254 1628 -213
rect 1521 -288 1556 -254
rect 1590 -288 1628 -254
rect 1521 -329 1628 -288
rect 1521 -363 1556 -329
rect 1590 -363 1628 -329
rect 1521 -404 1628 -363
rect 1521 -438 1556 -404
rect 1590 -438 1628 -404
rect 1521 -479 1628 -438
rect 1521 -513 1556 -479
rect 1590 -513 1628 -479
rect 1521 -554 1628 -513
rect 1521 -588 1556 -554
rect 1590 -588 1628 -554
rect 1521 -628 1628 -588
rect 1521 -662 1556 -628
rect 1590 -662 1628 -628
tri 1415 -674 1417 -672 sw
rect 1521 -674 1628 -662
rect 1731 64 1838 76
tri 1951 75 1952 76 ne
rect 1952 75 2061 76
tri 2061 75 2062 76 nw
tri 1952 74 1953 75 ne
rect 1731 30 1772 64
rect 1806 30 1838 64
rect 1731 -11 1838 30
rect 1731 -45 1772 -11
rect 1806 -45 1838 -11
rect 1731 -86 1838 -45
rect 1731 -120 1772 -86
rect 1806 -120 1838 -86
rect 1731 -161 1838 -120
rect 1731 -195 1772 -161
rect 1806 -195 1838 -161
rect 1731 -236 1838 -195
rect 1731 -270 1772 -236
rect 1806 -270 1838 -236
rect 1731 -311 1838 -270
rect 1731 -345 1772 -311
rect 1806 -345 1838 -311
rect 1731 -386 1838 -345
rect 1731 -420 1772 -386
rect 1806 -420 1838 -386
rect 1731 -461 1838 -420
rect 1731 -495 1772 -461
rect 1806 -495 1838 -461
rect 1731 -536 1838 -495
rect 1731 -570 1772 -536
rect 1806 -570 1838 -536
rect 1731 -611 1838 -570
rect 1731 -645 1772 -611
rect 1806 -645 1838 -611
tri 1729 -674 1731 -672 se
rect 1731 -674 1838 -645
rect 1953 46 2060 75
tri 2060 74 2061 75 nw
rect 1953 12 1988 46
rect 2022 12 2060 46
rect 1953 -29 2060 12
rect 1953 -63 1988 -29
rect 2022 -63 2060 -29
rect 1953 -104 2060 -63
rect 1953 -138 1988 -104
rect 2022 -138 2060 -104
rect 1953 -179 2060 -138
rect 1953 -213 1988 -179
rect 2022 -213 2060 -179
rect 1953 -254 2060 -213
rect 1953 -288 1988 -254
rect 2022 -288 2060 -254
rect 1953 -329 2060 -288
rect 1953 -363 1988 -329
rect 2022 -363 2060 -329
rect 1953 -404 2060 -363
rect 1953 -438 1988 -404
rect 2022 -438 2060 -404
rect 1953 -479 2060 -438
rect 1953 -513 1988 -479
rect 2022 -513 2060 -479
rect 1953 -554 2060 -513
rect 1953 -588 1988 -554
rect 2022 -588 2060 -554
rect 1953 -628 2060 -588
rect 1953 -662 1988 -628
rect 2022 -662 2060 -628
tri 1838 -674 1840 -672 sw
rect 1953 -674 2060 -662
rect 2163 64 2270 76
tri 2383 75 2384 76 ne
rect 2384 75 2493 76
tri 2493 75 2494 76 nw
tri 2384 74 2385 75 ne
rect 2163 30 2204 64
rect 2238 30 2270 64
rect 2163 -11 2270 30
rect 2163 -45 2204 -11
rect 2238 -45 2270 -11
rect 2163 -86 2270 -45
rect 2163 -120 2204 -86
rect 2238 -120 2270 -86
rect 2163 -161 2270 -120
rect 2163 -195 2204 -161
rect 2238 -195 2270 -161
rect 2163 -236 2270 -195
rect 2163 -270 2204 -236
rect 2238 -270 2270 -236
rect 2163 -311 2270 -270
rect 2163 -345 2204 -311
rect 2238 -345 2270 -311
rect 2163 -386 2270 -345
rect 2163 -420 2204 -386
rect 2238 -420 2270 -386
rect 2163 -461 2270 -420
rect 2163 -495 2204 -461
rect 2238 -495 2270 -461
rect 2163 -536 2270 -495
rect 2163 -570 2204 -536
rect 2238 -570 2270 -536
rect 2163 -611 2270 -570
rect 2163 -645 2204 -611
rect 2238 -645 2270 -611
tri 2161 -674 2163 -672 se
rect 2163 -674 2270 -645
rect 2385 46 2492 75
tri 2492 74 2493 75 nw
rect 2385 12 2420 46
rect 2454 12 2492 46
rect 2385 -29 2492 12
rect 2385 -63 2420 -29
rect 2454 -63 2492 -29
rect 2385 -104 2492 -63
rect 2385 -138 2420 -104
rect 2454 -138 2492 -104
rect 2385 -179 2492 -138
rect 2385 -213 2420 -179
rect 2454 -213 2492 -179
rect 2385 -254 2492 -213
rect 2385 -288 2420 -254
rect 2454 -288 2492 -254
rect 2385 -329 2492 -288
rect 2385 -363 2420 -329
rect 2454 -363 2492 -329
rect 2385 -404 2492 -363
rect 2385 -438 2420 -404
rect 2454 -438 2492 -404
rect 2385 -479 2492 -438
rect 2385 -513 2420 -479
rect 2454 -513 2492 -479
rect 2385 -554 2492 -513
rect 2385 -588 2420 -554
rect 2454 -588 2492 -554
rect 2385 -628 2492 -588
rect 2385 -662 2420 -628
rect 2454 -662 2492 -628
rect 2385 -674 2492 -662
rect 2630 64 2676 76
tri 2815 75 2816 76 ne
rect 2816 75 2925 76
tri 2925 75 2926 76 nw
tri 2816 74 2817 75 ne
rect 2630 30 2636 64
rect 2670 30 2676 64
rect 2630 -11 2676 30
rect 2630 -45 2636 -11
rect 2670 -45 2676 -11
rect 2630 -86 2676 -45
rect 2630 -120 2636 -86
rect 2670 -120 2676 -86
rect 2630 -161 2676 -120
rect 2630 -195 2636 -161
rect 2670 -195 2676 -161
rect 2630 -236 2676 -195
rect 2630 -270 2636 -236
rect 2670 -270 2676 -236
rect 2630 -311 2676 -270
rect 2630 -345 2636 -311
rect 2670 -345 2676 -311
rect 2630 -386 2676 -345
rect 2630 -420 2636 -386
rect 2670 -420 2676 -386
rect 2630 -461 2676 -420
rect 2630 -495 2636 -461
rect 2670 -495 2676 -461
rect 2630 -536 2676 -495
rect 2630 -570 2636 -536
rect 2670 -570 2676 -536
rect 2630 -611 2676 -570
rect 2630 -645 2636 -611
rect 2670 -645 2676 -611
rect 2630 -674 2676 -645
rect 2817 46 2924 75
tri 2924 74 2925 75 nw
rect 2817 12 2852 46
rect 2886 12 2924 46
rect 2817 -29 2924 12
rect 2817 -63 2852 -29
rect 2886 -63 2924 -29
rect 2817 -104 2924 -63
rect 2817 -138 2852 -104
rect 2886 -138 2924 -104
rect 2817 -179 2924 -138
rect 2817 -213 2852 -179
rect 2886 -213 2924 -179
rect 2817 -254 2924 -213
rect 2817 -288 2852 -254
rect 2886 -288 2924 -254
rect 2817 -329 2924 -288
rect 2817 -363 2852 -329
rect 2886 -363 2924 -329
rect 2817 -404 2924 -363
rect 2817 -438 2852 -404
rect 2886 -438 2924 -404
rect 2817 -479 2924 -438
rect 2817 -513 2852 -479
rect 2886 -513 2924 -479
rect 2817 -554 2924 -513
rect 2817 -588 2852 -554
rect 2886 -588 2924 -554
rect 2817 -628 2924 -588
rect 2817 -662 2852 -628
rect 2886 -662 2924 -628
tri 2676 -674 2678 -672 sw
rect 2817 -674 2924 -662
rect 3062 64 3108 76
tri 3276 75 3277 76 ne
rect 3277 75 3435 76
tri 3435 75 3436 76 nw
tri 3277 74 3278 75 ne
rect 3062 30 3068 64
rect 3102 30 3108 64
rect 3062 -11 3108 30
rect 3062 -45 3068 -11
rect 3102 -45 3108 -11
rect 3062 -86 3108 -45
rect 3062 -120 3068 -86
rect 3102 -120 3108 -86
rect 3062 -161 3108 -120
rect 3062 -195 3068 -161
rect 3102 -195 3108 -161
rect 3062 -236 3108 -195
rect 3062 -270 3068 -236
rect 3102 -270 3108 -236
rect 3062 -311 3108 -270
rect 3062 -345 3068 -311
rect 3102 -345 3108 -311
rect 3062 -386 3108 -345
rect 3062 -420 3068 -386
rect 3102 -420 3108 -386
rect 3062 -461 3108 -420
rect 3062 -495 3068 -461
rect 3102 -495 3108 -461
rect 3062 -536 3108 -495
rect 3062 -570 3068 -536
rect 3102 -570 3108 -536
rect 3062 -611 3108 -570
rect 3062 -645 3068 -611
rect 3102 -645 3108 -611
tri 3060 -674 3062 -672 se
rect 3062 -674 3108 -645
rect 3278 46 3434 75
tri 3434 74 3435 75 nw
rect 3278 12 3284 46
rect 3318 12 3394 46
rect 3428 12 3434 46
rect 3278 -29 3434 12
rect 3278 -63 3284 -29
rect 3318 -63 3394 -29
rect 3428 -63 3434 -29
rect 3278 -104 3434 -63
rect 3278 -138 3284 -104
rect 3318 -138 3394 -104
rect 3428 -138 3434 -104
rect 3278 -179 3434 -138
rect 3278 -213 3284 -179
rect 3318 -213 3394 -179
rect 3428 -213 3434 -179
rect 3278 -254 3434 -213
rect 3278 -288 3284 -254
rect 3318 -288 3394 -254
rect 3428 -288 3434 -254
rect 3278 -329 3434 -288
rect 3278 -363 3284 -329
rect 3318 -363 3394 -329
rect 3428 -363 3434 -329
rect 3278 -404 3434 -363
rect 3278 -438 3284 -404
rect 3318 -438 3394 -404
rect 3428 -438 3434 -404
rect 3278 -479 3434 -438
rect 3278 -513 3284 -479
rect 3318 -513 3394 -479
rect 3428 -513 3434 -479
rect 3278 -554 3434 -513
rect 3278 -588 3284 -554
rect 3318 -588 3394 -554
rect 3428 -588 3434 -554
rect 3278 -628 3434 -588
rect 3278 -662 3284 -628
rect 3318 -662 3394 -628
rect 3428 -662 3434 -628
rect 3278 -674 3434 -662
rect 3601 68 3760 76
rect 3653 16 3669 68
rect 3721 64 3760 68
rect 3754 30 3760 64
rect 3721 16 3760 30
rect 3601 1 3760 16
rect 3653 -51 3669 1
rect 3721 -11 3760 1
rect 3754 -45 3760 -11
rect 3721 -51 3760 -45
rect 3601 -66 3760 -51
rect 3653 -118 3669 -66
rect 3721 -86 3760 -66
rect 3601 -120 3610 -118
rect 3644 -120 3720 -118
rect 3754 -120 3760 -86
rect 3601 -133 3760 -120
rect 3653 -185 3669 -133
rect 3721 -161 3760 -133
rect 3601 -195 3610 -185
rect 3644 -195 3720 -185
rect 3754 -195 3760 -161
rect 3601 -200 3760 -195
rect 3653 -252 3669 -200
rect 3721 -236 3760 -200
rect 3601 -268 3610 -252
rect 3644 -268 3720 -252
rect 3653 -320 3669 -268
rect 3754 -270 3760 -236
rect 3721 -311 3760 -270
rect 3601 -336 3610 -320
rect 3644 -336 3720 -320
rect 3653 -388 3669 -336
rect 3754 -345 3760 -311
rect 3721 -386 3760 -345
rect 3601 -404 3610 -388
rect 3644 -404 3720 -388
rect 3653 -456 3669 -404
rect 3754 -420 3760 -386
rect 3721 -456 3760 -420
rect 3601 -461 3760 -456
rect 3601 -472 3610 -461
rect 3644 -472 3720 -461
rect 3653 -524 3669 -472
rect 3754 -495 3760 -461
rect 3721 -524 3760 -495
rect 3601 -536 3760 -524
rect 3601 -540 3610 -536
rect 3644 -540 3720 -536
rect 3653 -592 3669 -540
rect 3754 -570 3760 -536
rect 3721 -592 3760 -570
rect 3601 -608 3760 -592
rect 3653 -660 3669 -608
rect 3721 -611 3760 -608
rect 3754 -645 3760 -611
rect 3721 -660 3760 -645
rect 38 -677 86 -674
tri 86 -677 89 -674 sw
tri 439 -677 442 -674 se
rect 442 -677 553 -674
tri 553 -677 556 -674 sw
tri 806 -677 809 -674 se
rect 809 -677 956 -674
rect 38 -684 89 -677
tri 89 -684 96 -677 sw
tri 432 -684 439 -677 se
rect 439 -684 556 -677
tri 556 -684 563 -677 sw
tri 799 -684 806 -677 se
rect 806 -684 956 -677
rect 38 -686 96 -684
tri 96 -686 98 -684 sw
tri 430 -686 432 -684 se
rect 432 -686 563 -684
tri 563 -686 565 -684 sw
tri 797 -686 799 -684 se
rect 799 -686 956 -684
rect 38 -687 98 -686
rect 38 -721 44 -687
rect 78 -706 98 -687
tri 98 -706 118 -686 sw
tri 410 -706 430 -686 se
rect 430 -706 476 -686
rect 78 -720 476 -706
rect 510 -706 565 -686
tri 565 -706 585 -686 sw
tri 777 -706 797 -686 se
rect 797 -706 908 -686
rect 510 -720 908 -706
rect 942 -720 956 -686
rect 1308 -677 1417 -674
tri 1417 -677 1420 -674 sw
tri 1726 -677 1729 -674 se
rect 1729 -677 1840 -674
tri 1840 -677 1843 -674 sw
tri 2158 -677 2161 -674 se
rect 2161 -677 2270 -674
rect 1308 -684 1420 -677
tri 1420 -684 1427 -677 sw
tri 1719 -684 1726 -677 se
rect 1726 -684 1843 -677
tri 1843 -684 1850 -677 sw
tri 2151 -684 2158 -677 se
rect 2158 -684 2270 -677
rect 1308 -686 1427 -684
tri 1427 -686 1429 -684 sw
tri 1717 -686 1719 -684 se
rect 1719 -686 1850 -684
tri 1850 -686 1852 -684 sw
tri 2149 -686 2151 -684 se
rect 2151 -686 2270 -684
tri 1297 -706 1308 -695 se
rect 1308 -706 1340 -686
tri 1283 -720 1297 -706 se
rect 1297 -720 1340 -706
rect 1374 -706 1429 -686
tri 1429 -706 1449 -686 sw
tri 1697 -706 1717 -686 se
rect 1717 -706 1772 -686
rect 1374 -720 1772 -706
rect 1806 -698 1852 -686
tri 1852 -698 1864 -686 sw
tri 2137 -698 2149 -686 se
rect 2149 -698 2204 -686
rect 1806 -706 1864 -698
tri 1864 -706 1872 -698 sw
tri 2129 -706 2137 -698 se
rect 2137 -706 2204 -698
rect 1806 -720 2204 -706
rect 2238 -706 2270 -686
rect 2630 -677 2678 -674
tri 2678 -677 2681 -674 sw
tri 3057 -677 3060 -674 se
rect 3060 -677 3108 -674
rect 2630 -684 2681 -677
tri 2681 -684 2688 -677 sw
tri 3050 -684 3057 -677 se
rect 3057 -684 3108 -677
rect 2630 -686 2688 -684
tri 2688 -686 2690 -684 sw
tri 3048 -686 3050 -684 se
rect 3050 -686 3108 -684
tri 2270 -706 2281 -695 sw
rect 2238 -720 2281 -706
tri 2281 -720 2295 -706 sw
rect 2630 -720 2636 -686
rect 2670 -706 2690 -686
tri 2690 -706 2710 -686 sw
tri 3028 -706 3048 -686 se
rect 3048 -706 3068 -686
rect 2670 -720 3068 -706
rect 3102 -720 3108 -686
rect 78 -721 956 -720
rect 38 -760 956 -721
tri 1243 -760 1283 -720 se
rect 1283 -760 2295 -720
tri 2295 -760 2335 -720 sw
rect 2630 -730 3108 -720
rect 3601 -676 3760 -660
rect 38 -794 44 -760
rect 78 -794 476 -760
rect 510 -794 908 -760
rect 942 -794 956 -760
tri 1209 -794 1243 -760 se
rect 1243 -794 1340 -760
rect 1374 -794 1772 -760
rect 1806 -794 2204 -760
rect 2238 -794 2335 -760
tri 2335 -794 2369 -760 sw
rect 2630 -794 2636 -730
rect 2688 -782 2700 -730
rect 2752 -760 3108 -730
tri 3567 -757 3601 -723 se
rect 3653 -728 3669 -676
rect 3721 -686 3760 -676
rect 3754 -720 3760 -686
rect 3721 -728 3760 -720
rect 3927 70 4086 76
rect 3979 64 4086 70
rect 3979 30 4046 64
rect 4080 30 4086 64
rect 3979 18 4086 30
rect 3927 6 4086 18
rect 3979 -11 4086 6
rect 3979 -45 4046 -11
rect 4080 -45 4086 -11
rect 3979 -46 4086 -45
rect 3927 -86 4086 -46
rect 3927 -120 3936 -86
rect 3970 -120 4046 -86
rect 4080 -120 4086 -86
rect 3927 -161 4086 -120
rect 3927 -195 3936 -161
rect 3970 -195 4046 -161
rect 4080 -195 4086 -161
rect 3927 -236 4086 -195
rect 3927 -270 3936 -236
rect 3970 -270 4046 -236
rect 4080 -270 4086 -236
rect 3927 -311 4086 -270
rect 3927 -345 3936 -311
rect 3970 -345 4046 -311
rect 4080 -345 4086 -311
rect 3927 -386 4086 -345
rect 3927 -420 3936 -386
rect 3970 -420 4046 -386
rect 4080 -420 4086 -386
rect 3927 -461 4086 -420
rect 3927 -495 3936 -461
rect 3970 -495 4046 -461
rect 4080 -495 4086 -461
rect 3927 -536 4086 -495
rect 3927 -570 3936 -536
rect 3970 -570 4046 -536
rect 4080 -570 4086 -536
rect 3927 -611 4086 -570
rect 3927 -645 3936 -611
rect 3970 -645 4046 -611
rect 4080 -645 4086 -611
rect 3927 -686 4086 -645
rect 3927 -720 3936 -686
rect 3970 -720 4046 -686
rect 4080 -720 4086 -686
rect 3601 -744 3760 -728
tri 3564 -760 3567 -757 se
rect 3567 -760 3601 -757
rect 2752 -782 3068 -760
rect 2670 -794 3068 -782
rect 3102 -794 3108 -760
tri 3530 -794 3564 -760 se
rect 3564 -794 3601 -760
rect 38 -806 956 -794
tri 1197 -806 1209 -794 se
rect 1209 -806 2369 -794
tri 2369 -806 2381 -794 sw
rect 2630 -806 3108 -794
tri 3518 -806 3530 -794 se
rect 3530 -796 3601 -794
rect 3653 -796 3669 -744
rect 3721 -757 3760 -744
tri 3760 -757 3794 -723 sw
tri 3893 -757 3927 -723 se
rect 3927 -757 4086 -720
rect 4253 70 4305 76
rect 4253 6 4305 18
rect 4540 -2 4546 50
rect 4598 -2 4610 50
rect 4662 41 5102 50
rect 4662 7 4984 41
rect 5018 7 5056 41
rect 5090 7 5102 41
rect 4662 -2 5102 7
rect 5356 19 5402 108
tri 5402 100 5410 108 nw
rect 5666 89 5675 109
rect 5709 89 5718 109
rect 5666 33 5718 37
rect 5356 -15 5362 19
rect 5396 -15 5402 19
rect 4253 -86 4305 -46
rect 5265 -38 5317 -32
rect 4253 -120 4262 -86
rect 4296 -120 4305 -86
tri 5255 -90 5265 -80 se
tri 5253 -92 5255 -90 se
rect 5255 -92 5317 -90
tri 5235 -110 5253 -92 se
rect 5253 -102 5317 -92
rect 5253 -110 5265 -102
rect 4253 -161 4305 -120
rect 4253 -195 4262 -161
rect 4296 -195 4305 -161
rect 4459 -163 4465 -111
rect 4517 -163 4529 -111
rect 4581 -163 4589 -111
rect 4673 -119 4807 -110
rect 4859 -119 4871 -110
rect 4673 -153 4685 -119
rect 4719 -153 4777 -119
rect 4859 -153 4868 -119
rect 4673 -162 4807 -153
rect 4859 -162 4871 -153
rect 4923 -162 4929 -110
tri 5231 -114 5235 -110 se
rect 5235 -114 5265 -110
rect 4985 -120 5265 -114
rect 4985 -154 4997 -120
rect 5031 -154 5081 -120
rect 5115 -154 5165 -120
rect 5199 -154 5265 -120
rect 4985 -160 5317 -154
rect 5356 -56 5402 -15
rect 5356 -90 5362 -56
rect 5396 -90 5402 -56
rect 5356 -131 5402 -90
rect 4253 -236 4305 -195
rect 5356 -165 5362 -131
rect 5396 -165 5402 -131
rect 5356 -206 5402 -165
tri 5214 -236 5244 -206 se
rect 5244 -212 5296 -206
rect 4253 -270 4262 -236
rect 4296 -270 4305 -236
rect 4253 -311 4305 -270
rect 4253 -345 4262 -311
rect 4296 -345 4305 -311
rect 4253 -386 4305 -345
rect 4253 -420 4262 -386
rect 4296 -420 4305 -386
rect 4253 -461 4305 -420
rect 4253 -495 4262 -461
rect 4296 -495 4305 -461
rect 4253 -536 4305 -495
rect 4253 -570 4262 -536
rect 4296 -570 4305 -536
rect 4253 -611 4305 -570
rect 4253 -645 4262 -611
rect 4296 -645 4305 -611
rect 4253 -686 4305 -645
rect 4253 -720 4262 -686
rect 4296 -720 4305 -686
rect 4363 -258 4415 -252
rect 4363 -322 4415 -310
rect 4778 -264 5244 -236
rect 4778 -276 5296 -264
rect 4778 -310 4784 -276
rect 4818 -310 5096 -276
rect 5130 -310 5244 -276
rect 4778 -328 5244 -310
rect 4778 -334 5296 -328
rect 5356 -240 5362 -206
rect 5396 -240 5402 -206
rect 5356 -281 5402 -240
rect 5356 -315 5362 -281
rect 5396 -315 5402 -281
rect 4778 -351 4841 -334
tri 4841 -351 4858 -334 nw
tri 5056 -351 5073 -334 ne
rect 5073 -351 5153 -334
tri 5153 -351 5170 -334 nw
rect 4363 -415 4415 -374
rect 4363 -449 4372 -415
rect 4406 -449 4415 -415
rect 4363 -491 4415 -449
rect 4363 -525 4372 -491
rect 4406 -525 4415 -491
rect 4363 -567 4415 -525
rect 4363 -601 4372 -567
rect 4406 -601 4415 -567
rect 4363 -643 4415 -601
rect 4363 -677 4372 -643
rect 4406 -677 4415 -643
rect 4363 -689 4415 -677
rect 4622 -381 4668 -369
rect 4622 -415 4628 -381
rect 4662 -415 4668 -381
rect 4622 -456 4668 -415
rect 4622 -490 4628 -456
rect 4662 -490 4668 -456
rect 4622 -532 4668 -490
rect 4622 -566 4628 -532
rect 4662 -566 4668 -532
rect 4622 -608 4668 -566
rect 4622 -642 4628 -608
rect 4662 -642 4668 -608
rect 4622 -684 4668 -642
tri 4086 -757 4120 -723 sw
tri 4219 -757 4253 -723 se
rect 4253 -757 4305 -720
rect 4622 -718 4628 -684
rect 4662 -718 4668 -684
rect 4778 -385 4784 -351
rect 4818 -385 4824 -351
tri 4824 -368 4841 -351 nw
tri 5073 -368 5090 -351 ne
rect 4778 -427 4824 -385
rect 4778 -461 4784 -427
rect 4818 -461 4824 -427
rect 4778 -503 4824 -461
rect 4778 -537 4784 -503
rect 4818 -537 4824 -503
rect 4778 -579 4824 -537
rect 4778 -613 4784 -579
rect 4818 -613 4824 -579
rect 4778 -655 4824 -613
rect 4778 -689 4784 -655
rect 4818 -689 4824 -655
rect 4778 -701 4824 -689
rect 4934 -381 4980 -369
rect 4934 -415 4940 -381
rect 4974 -415 4980 -381
rect 4934 -456 4980 -415
rect 4934 -490 4940 -456
rect 4974 -490 4980 -456
rect 4934 -532 4980 -490
rect 4934 -566 4940 -532
rect 4974 -566 4980 -532
rect 4934 -608 4980 -566
rect 4934 -642 4940 -608
rect 4974 -642 4980 -608
rect 4934 -684 4980 -642
tri 4305 -757 4339 -723 sw
tri 4588 -757 4622 -723 se
rect 4622 -757 4668 -718
rect 4934 -718 4940 -684
rect 4974 -718 4980 -684
rect 5090 -385 5096 -351
rect 5130 -356 5148 -351
tri 5148 -356 5153 -351 nw
rect 5356 -356 5402 -315
rect 5130 -385 5136 -356
tri 5136 -368 5148 -356 nw
rect 5090 -427 5136 -385
rect 5090 -461 5096 -427
rect 5130 -461 5136 -427
rect 5090 -503 5136 -461
rect 5090 -537 5096 -503
rect 5130 -537 5136 -503
rect 5090 -579 5136 -537
rect 5090 -613 5096 -579
rect 5130 -613 5136 -579
rect 5090 -655 5136 -613
rect 5090 -689 5096 -655
rect 5130 -689 5136 -655
rect 5090 -701 5136 -689
rect 5246 -381 5292 -369
rect 5246 -415 5252 -381
rect 5286 -415 5292 -381
rect 5246 -456 5292 -415
rect 5246 -490 5252 -456
rect 5286 -490 5292 -456
rect 5246 -532 5292 -490
rect 5246 -566 5252 -532
rect 5286 -566 5292 -532
rect 5246 -608 5292 -566
rect 5246 -642 5252 -608
rect 5286 -642 5292 -608
rect 5356 -390 5362 -356
rect 5396 -390 5402 -356
rect 5356 -431 5402 -390
rect 5356 -465 5362 -431
rect 5396 -465 5402 -431
rect 5356 -506 5402 -465
rect 5356 -540 5362 -506
rect 5396 -540 5402 -506
rect 5356 -582 5402 -540
rect 5356 -616 5362 -582
rect 5396 -616 5402 -582
rect 5356 -628 5402 -616
rect 5512 19 5558 31
rect 5512 -15 5518 19
rect 5552 -15 5558 19
rect 5512 -58 5558 -15
rect 5512 -92 5518 -58
rect 5552 -92 5558 -58
rect 5512 -136 5558 -92
rect 5512 -170 5518 -136
rect 5552 -170 5558 -136
rect 5512 -214 5558 -170
rect 5512 -248 5518 -214
rect 5552 -248 5558 -214
rect 5512 -292 5558 -248
rect 5512 -326 5518 -292
rect 5552 -326 5558 -292
rect 5512 -370 5558 -326
rect 5512 -404 5518 -370
rect 5552 -404 5558 -370
rect 5512 -448 5558 -404
rect 5512 -482 5518 -448
rect 5552 -482 5558 -448
rect 5512 -526 5558 -482
rect 5512 -560 5518 -526
rect 5552 -560 5558 -526
rect 5512 -604 5558 -560
rect 5246 -684 5292 -642
tri 4668 -757 4702 -723 sw
tri 4900 -757 4934 -723 se
rect 4934 -757 4980 -718
rect 5246 -718 5252 -684
rect 5286 -718 5292 -684
tri 4980 -757 5014 -723 sw
tri 5212 -757 5246 -723 se
rect 5246 -757 5292 -718
rect 5512 -638 5518 -604
rect 5552 -638 5558 -604
rect 5666 25 5675 33
rect 5709 25 5718 33
rect 5666 -43 5718 -27
rect 5666 -77 5675 -43
rect 5709 -77 5718 -43
rect 5666 -120 5718 -77
rect 5666 -154 5675 -120
rect 5709 -154 5718 -120
rect 5666 -197 5718 -154
rect 5666 -231 5675 -197
rect 5709 -231 5718 -197
rect 5666 -274 5718 -231
rect 5666 -308 5675 -274
rect 5709 -308 5718 -274
rect 5666 -351 5718 -308
rect 5666 -385 5675 -351
rect 5709 -385 5718 -351
rect 5666 -428 5718 -385
rect 5666 -462 5675 -428
rect 5709 -462 5718 -428
rect 5666 -505 5718 -462
rect 5666 -539 5675 -505
rect 5709 -539 5718 -505
rect 5666 -582 5718 -539
rect 5666 -616 5675 -582
rect 5709 -616 5718 -582
rect 5666 -628 5718 -616
rect 5512 -682 5558 -638
rect 5512 -716 5518 -682
rect 5552 -716 5558 -682
tri 5292 -757 5326 -723 sw
tri 5478 -757 5512 -723 se
rect 5512 -757 5558 -716
tri 5558 -757 5592 -723 sw
rect 3721 -760 5752 -757
rect 3754 -794 3936 -760
rect 3970 -794 4046 -760
rect 4080 -794 4262 -760
rect 4296 -794 4628 -760
rect 4662 -794 4940 -760
rect 4974 -794 5252 -760
rect 5286 -794 5518 -760
rect 5552 -794 5752 -760
rect 3721 -796 5752 -794
rect 3530 -806 5752 -796
tri 1131 -872 1197 -806 se
rect 1197 -838 2381 -806
tri 2381 -838 2413 -806 sw
tri 3486 -838 3518 -806 se
rect 3518 -812 5752 -806
rect 3518 -838 3601 -812
rect 1197 -872 2413 -838
tri 2413 -872 2447 -838 sw
tri 3452 -872 3486 -838 se
rect 3486 -864 3601 -838
rect 3653 -864 3669 -812
rect 3721 -864 5752 -812
rect 3486 -872 5752 -864
rect 14 -878 5752 -872
rect 14 -912 67 -878
rect 101 -912 140 -878
rect 174 -912 213 -878
rect 247 -912 286 -878
rect 320 -912 359 -878
rect 393 -912 432 -878
rect 466 -912 505 -878
rect 539 -912 578 -878
rect 612 -912 651 -878
rect 685 -912 724 -878
rect 758 -912 797 -878
rect 831 -912 870 -878
rect 904 -912 943 -878
rect 977 -912 1016 -878
rect 1050 -912 1089 -878
rect 1123 -912 1162 -878
rect 1196 -912 1235 -878
rect 1269 -912 1308 -878
rect 1342 -912 1381 -878
rect 1415 -912 1454 -878
rect 1488 -912 1527 -878
rect 1561 -912 1600 -878
rect 1634 -912 1673 -878
rect 1707 -912 1746 -878
rect 1780 -912 1819 -878
rect 1853 -912 1892 -878
rect 1926 -912 1965 -878
rect 1999 -912 2038 -878
rect 2072 -912 2111 -878
rect 2145 -912 2184 -878
rect 2218 -912 2257 -878
rect 2291 -912 2330 -878
rect 2364 -912 2403 -878
rect 2437 -912 2476 -878
rect 2510 -912 2549 -878
rect 2583 -912 2622 -878
rect 2656 -912 2695 -878
rect 2729 -912 2768 -878
rect 2802 -912 2841 -878
rect 2875 -912 2914 -878
rect 2948 -912 2987 -878
rect 3021 -912 3060 -878
rect 3094 -912 3133 -878
rect 3167 -912 3206 -878
rect 3240 -912 3279 -878
rect 3313 -912 3352 -878
rect 3386 -912 3425 -878
rect 3459 -912 3498 -878
rect 3532 -912 3570 -878
rect 3604 -880 3642 -878
rect 3676 -880 3714 -878
rect 3748 -912 3786 -878
rect 3820 -912 3858 -878
rect 3892 -912 3930 -878
rect 3964 -912 4002 -878
rect 4036 -912 4074 -878
rect 4108 -912 4146 -878
rect 4180 -912 4218 -878
rect 4252 -912 4290 -878
rect 4324 -912 4362 -878
rect 4396 -912 4434 -878
rect 4468 -912 4506 -878
rect 4540 -912 4578 -878
rect 4612 -912 4650 -878
rect 4684 -912 4722 -878
rect 4756 -912 4794 -878
rect 4828 -912 4866 -878
rect 4900 -912 4938 -878
rect 4972 -912 5010 -878
rect 5044 -912 5082 -878
rect 5116 -912 5154 -878
rect 5188 -912 5226 -878
rect 5260 -912 5298 -878
rect 5332 -912 5370 -878
rect 5404 -912 5442 -878
rect 5476 -912 5514 -878
rect 5548 -912 5586 -878
rect 5620 -912 5658 -878
rect 5692 -912 5752 -878
rect 14 -932 3601 -912
rect 3653 -932 3669 -912
rect 3721 -932 5752 -912
rect 14 -1172 5752 -932
<< via1 >>
rect 703 2135 755 2173
rect 703 2121 712 2135
rect 712 2121 746 2135
rect 746 2121 755 2135
rect 703 2059 755 2091
rect 703 2039 712 2059
rect 712 2039 746 2059
rect 746 2039 755 2059
rect 703 1983 755 2008
rect 703 1956 712 1983
rect 712 1956 746 1983
rect 746 1956 755 1983
rect 703 1907 755 1925
rect 703 1873 712 1907
rect 712 1873 746 1907
rect 746 1873 755 1907
rect 1763 2135 1815 2166
rect 1763 2114 1772 2135
rect 1772 2114 1806 2135
rect 1806 2114 1815 2135
rect 1763 2059 1815 2084
rect 1763 2032 1772 2059
rect 1772 2032 1806 2059
rect 1806 2032 1815 2059
rect 1763 1983 1815 2002
rect 1763 1950 1772 1983
rect 1772 1950 1806 1983
rect 1806 1950 1815 1983
rect 1763 1907 1815 1919
rect 1763 1873 1772 1907
rect 1772 1873 1806 1907
rect 1806 1873 1815 1907
rect 1763 1867 1815 1873
rect 2075 2135 2127 2166
rect 2075 2114 2084 2135
rect 2084 2114 2118 2135
rect 2118 2114 2127 2135
rect 2075 2059 2127 2084
rect 2075 2032 2084 2059
rect 2084 2032 2118 2059
rect 2118 2032 2127 2059
rect 2075 1983 2127 2002
rect 2075 1950 2084 1983
rect 2084 1950 2118 1983
rect 2118 1950 2127 1983
rect 2075 1907 2127 1919
rect 2075 1873 2084 1907
rect 2084 1873 2118 1907
rect 2118 1873 2127 1907
rect 2075 1867 2127 1873
rect 3637 2359 3689 2365
rect 3637 2325 3646 2359
rect 3646 2325 3680 2359
rect 3680 2325 3689 2359
rect 3637 2313 3689 2325
rect 3392 2296 3444 2305
rect 3392 2262 3396 2296
rect 3396 2262 3430 2296
rect 3430 2262 3444 2296
rect 3392 2253 3444 2262
rect 3456 2296 3508 2305
rect 3456 2262 3468 2296
rect 3468 2262 3502 2296
rect 3502 2262 3508 2296
rect 3456 2253 3508 2262
rect 3637 2287 3689 2301
rect 3637 2253 3646 2287
rect 3646 2253 3680 2287
rect 3680 2253 3689 2287
rect 3885 2358 3937 2364
rect 3885 2324 3894 2358
rect 3894 2324 3928 2358
rect 3928 2324 3937 2358
rect 3885 2312 3937 2324
rect 3885 2286 3937 2300
rect 3637 2249 3689 2253
rect 3885 2252 3894 2286
rect 3894 2252 3928 2286
rect 3928 2252 3937 2286
rect 3885 2248 3937 2252
rect 3601 2102 3653 2154
rect 3669 2102 3721 2154
rect 3601 2027 3653 2079
rect 3669 2027 3721 2079
rect 3601 1951 3653 2003
rect 3669 1951 3721 2003
rect 131 1817 183 1825
rect 131 1783 137 1817
rect 137 1783 171 1817
rect 171 1783 183 1817
rect 131 1773 183 1783
rect 195 1817 247 1825
rect 195 1783 231 1817
rect 231 1783 247 1817
rect 195 1773 247 1783
rect 549 1817 601 1826
rect 613 1817 665 1826
rect 549 1783 578 1817
rect 578 1783 601 1817
rect 613 1783 650 1817
rect 650 1783 665 1817
rect 549 1774 601 1783
rect 613 1774 665 1783
rect 1042 1817 1094 1826
rect 1106 1817 1158 1826
rect 1042 1783 1084 1817
rect 1084 1783 1094 1817
rect 1106 1783 1118 1817
rect 1118 1783 1158 1817
rect 1042 1774 1094 1783
rect 1106 1774 1158 1783
rect 1563 1773 1615 1825
rect 1627 1817 1679 1825
rect 1627 1783 1673 1817
rect 1673 1783 1679 1817
rect 1627 1773 1679 1783
rect 2290 1817 2342 1825
rect 2290 1783 2306 1817
rect 2306 1783 2340 1817
rect 2340 1783 2342 1817
rect 2290 1773 2342 1783
rect 2354 1817 2406 1825
rect 2354 1783 2378 1817
rect 2378 1783 2406 1817
rect 2354 1773 2406 1783
rect 2506 1817 2558 1826
rect 2506 1783 2510 1817
rect 2510 1783 2544 1817
rect 2544 1783 2558 1817
rect 2506 1774 2558 1783
rect 2570 1817 2622 1826
rect 2570 1783 2582 1817
rect 2582 1783 2616 1817
rect 2616 1783 2622 1817
rect 2570 1774 2622 1783
rect 2791 1817 2843 1826
rect 2791 1783 2795 1817
rect 2795 1783 2829 1817
rect 2829 1783 2843 1817
rect 2791 1774 2843 1783
rect 2855 1817 2907 1826
rect 2855 1783 2867 1817
rect 2867 1783 2901 1817
rect 2901 1783 2907 1817
rect 2855 1774 2907 1783
rect 2981 1817 3033 1826
rect 2981 1783 2987 1817
rect 2987 1783 3021 1817
rect 3021 1783 3033 1817
rect 2981 1774 3033 1783
rect 3045 1817 3097 1826
rect 3045 1783 3059 1817
rect 3059 1783 3093 1817
rect 3093 1783 3097 1817
rect 3045 1774 3097 1783
rect 3236 1790 3288 1842
rect 3300 1790 3352 1842
rect 131 1673 183 1725
rect 195 1673 247 1725
rect 2290 1673 2342 1725
rect 2354 1673 2406 1725
rect 3392 1673 3444 1725
rect 3456 1673 3508 1725
rect 4883 1673 4935 1725
rect 4947 1673 4999 1725
rect 1042 1513 1094 1565
rect 1106 1513 1158 1565
rect 1563 1513 1615 1565
rect 1627 1513 1679 1565
rect 3891 1513 3943 1565
rect 3955 1513 4007 1565
rect 1192 1433 1244 1485
rect 1256 1433 1308 1485
rect 4293 1433 4345 1485
rect 4357 1433 4409 1485
rect 709 1353 761 1405
rect 773 1353 825 1405
rect 2506 1353 2558 1405
rect 2570 1353 2622 1405
rect 2728 1353 2780 1405
rect 2792 1353 2844 1405
rect 4576 1353 4628 1405
rect 4640 1353 4692 1405
rect 1719 1273 1771 1325
rect 1783 1273 1835 1325
rect 2594 1273 2646 1325
rect 2658 1273 2710 1325
rect 2081 1193 2133 1245
rect 2145 1193 2197 1245
rect 4470 1193 4522 1245
rect 4534 1193 4586 1245
rect 3767 1109 3819 1161
rect 3831 1109 3883 1161
rect 3236 796 3288 848
rect 3300 796 3352 848
rect 5636 796 5688 848
rect 5700 796 5752 848
rect 2981 678 3033 730
rect 3045 678 3097 730
rect 5480 678 5532 730
rect 5544 678 5596 730
rect 2878 592 2930 644
rect 5377 598 5429 650
rect 5441 598 5493 650
rect 2878 528 2930 580
rect 4459 495 4511 547
rect 4459 431 4511 483
rect 549 333 601 385
rect 613 333 665 385
rect 1875 333 1927 385
rect 1939 333 1991 385
rect 549 280 601 289
rect 613 280 665 289
rect 549 246 574 280
rect 574 246 601 280
rect 613 246 651 280
rect 651 246 665 280
rect 549 237 601 246
rect 613 237 665 246
rect 1192 280 1244 289
rect 1192 246 1198 280
rect 1198 246 1232 280
rect 1232 246 1244 280
rect 1192 237 1244 246
rect 1258 280 1310 289
rect 1258 246 1270 280
rect 1270 246 1304 280
rect 1304 246 1310 280
rect 1258 237 1310 246
rect 1875 280 1927 289
rect 1875 246 1877 280
rect 1877 246 1911 280
rect 1911 246 1927 280
rect 1875 237 1927 246
rect 1939 280 1991 289
rect 1939 246 1954 280
rect 1954 246 1988 280
rect 1988 246 1991 280
rect 1939 237 1991 246
rect 2804 280 2856 289
rect 2804 246 2819 280
rect 2819 246 2853 280
rect 2853 246 2856 280
rect 2804 237 2856 246
rect 2868 280 2920 289
rect 2868 246 2896 280
rect 2896 246 2920 280
rect 2868 237 2920 246
rect 3795 280 3847 289
rect 3795 246 3799 280
rect 3799 246 3833 280
rect 3833 246 3847 280
rect 3795 237 3847 246
rect 3859 280 3911 289
rect 3859 246 3871 280
rect 3871 246 3905 280
rect 3905 246 3911 280
rect 3859 237 3911 246
rect 4183 280 4235 289
rect 4183 246 4197 280
rect 4197 246 4231 280
rect 4231 246 4235 280
rect 4183 237 4235 246
rect 4247 237 4299 289
rect 4652 285 4704 289
rect 4716 285 4768 289
rect 4652 251 4669 285
rect 4669 251 4704 285
rect 4716 251 4742 285
rect 4742 251 4768 285
rect 4652 237 4704 251
rect 4716 237 4768 251
rect 5195 239 5247 291
rect 5259 239 5311 291
rect 5377 280 5429 292
rect 5441 280 5493 292
rect 5377 246 5394 280
rect 5394 246 5429 280
rect 5441 246 5467 280
rect 5467 246 5493 280
rect 5377 240 5429 246
rect 5441 240 5493 246
rect 5556 280 5608 289
rect 5620 280 5672 289
rect 5556 246 5577 280
rect 5577 246 5608 280
rect 5620 246 5649 280
rect 5649 246 5672 280
rect 5556 237 5608 246
rect 5620 237 5672 246
rect -461 -638 -409 -586
rect -376 -638 -324 -586
rect -291 -638 -239 -586
rect -207 -638 -155 -586
rect -123 -638 -71 -586
rect -461 -748 -409 -696
rect -376 -748 -324 -696
rect -291 -748 -239 -696
rect -207 -748 -155 -696
rect -123 -748 -71 -696
rect 827 18 879 70
rect 903 64 955 70
rect 903 30 908 64
rect 908 30 942 64
rect 942 30 955 64
rect 903 18 955 30
rect 827 -71 879 -19
rect 903 -45 908 -19
rect 908 -45 942 -19
rect 942 -45 955 -19
rect 903 -71 955 -45
rect 827 -160 879 -108
rect 903 -120 908 -108
rect 908 -120 942 -108
rect 942 -120 955 -108
rect 903 -160 955 -120
rect 827 -249 879 -197
rect 903 -236 955 -197
rect 903 -249 908 -236
rect 908 -249 942 -236
rect 942 -249 955 -236
rect 3601 64 3653 68
rect 3601 30 3610 64
rect 3610 30 3644 64
rect 3644 30 3653 64
rect 3601 16 3653 30
rect 3669 64 3721 68
rect 3669 30 3720 64
rect 3720 30 3721 64
rect 3669 16 3721 30
rect 3601 -11 3653 1
rect 3601 -45 3610 -11
rect 3610 -45 3644 -11
rect 3644 -45 3653 -11
rect 3601 -51 3653 -45
rect 3669 -11 3721 1
rect 3669 -45 3720 -11
rect 3720 -45 3721 -11
rect 3669 -51 3721 -45
rect 3601 -86 3653 -66
rect 3601 -118 3610 -86
rect 3610 -118 3644 -86
rect 3644 -118 3653 -86
rect 3669 -86 3721 -66
rect 3669 -118 3720 -86
rect 3720 -118 3721 -86
rect 3601 -161 3653 -133
rect 3601 -185 3610 -161
rect 3610 -185 3644 -161
rect 3644 -185 3653 -161
rect 3669 -161 3721 -133
rect 3669 -185 3720 -161
rect 3720 -185 3721 -161
rect 3601 -236 3653 -200
rect 3601 -252 3610 -236
rect 3610 -252 3644 -236
rect 3644 -252 3653 -236
rect 3669 -236 3721 -200
rect 3669 -252 3720 -236
rect 3720 -252 3721 -236
rect 3601 -270 3610 -268
rect 3610 -270 3644 -268
rect 3644 -270 3653 -268
rect 3601 -311 3653 -270
rect 3601 -320 3610 -311
rect 3610 -320 3644 -311
rect 3644 -320 3653 -311
rect 3669 -270 3720 -268
rect 3720 -270 3721 -268
rect 3669 -311 3721 -270
rect 3669 -320 3720 -311
rect 3720 -320 3721 -311
rect 3601 -345 3610 -336
rect 3610 -345 3644 -336
rect 3644 -345 3653 -336
rect 3601 -386 3653 -345
rect 3601 -388 3610 -386
rect 3610 -388 3644 -386
rect 3644 -388 3653 -386
rect 3669 -345 3720 -336
rect 3720 -345 3721 -336
rect 3669 -386 3721 -345
rect 3669 -388 3720 -386
rect 3720 -388 3721 -386
rect 3601 -420 3610 -404
rect 3610 -420 3644 -404
rect 3644 -420 3653 -404
rect 3601 -456 3653 -420
rect 3669 -420 3720 -404
rect 3720 -420 3721 -404
rect 3669 -456 3721 -420
rect 3601 -495 3610 -472
rect 3610 -495 3644 -472
rect 3644 -495 3653 -472
rect 3601 -524 3653 -495
rect 3669 -495 3720 -472
rect 3720 -495 3721 -472
rect 3669 -524 3721 -495
rect 3601 -570 3610 -540
rect 3610 -570 3644 -540
rect 3644 -570 3653 -540
rect 3601 -592 3653 -570
rect 3669 -570 3720 -540
rect 3720 -570 3721 -540
rect 3669 -592 3721 -570
rect 3601 -611 3653 -608
rect 3601 -645 3610 -611
rect 3610 -645 3644 -611
rect 3644 -645 3653 -611
rect 3601 -660 3653 -645
rect 3669 -611 3721 -608
rect 3669 -645 3720 -611
rect 3720 -645 3721 -611
rect 3669 -660 3721 -645
rect 3601 -686 3653 -676
rect 3601 -720 3610 -686
rect 3610 -720 3644 -686
rect 3644 -720 3653 -686
rect 2636 -760 2688 -730
rect 2636 -782 2670 -760
rect 2670 -782 2688 -760
rect 2700 -782 2752 -730
rect 3601 -728 3653 -720
rect 3669 -686 3721 -676
rect 3669 -720 3720 -686
rect 3720 -720 3721 -686
rect 3669 -728 3721 -720
rect 3927 64 3979 70
rect 3927 30 3936 64
rect 3936 30 3970 64
rect 3970 30 3979 64
rect 3927 18 3979 30
rect 3927 -11 3979 6
rect 3927 -45 3936 -11
rect 3936 -45 3970 -11
rect 3970 -45 3979 -11
rect 3927 -46 3979 -45
rect 3601 -760 3653 -744
rect 3601 -794 3610 -760
rect 3610 -794 3644 -760
rect 3644 -794 3653 -760
rect 3601 -796 3653 -794
rect 3669 -760 3721 -744
rect 4253 64 4305 70
rect 4253 30 4262 64
rect 4262 30 4296 64
rect 4296 30 4305 64
rect 4253 18 4305 30
rect 4253 -11 4305 6
rect 4546 41 4598 50
rect 4546 7 4552 41
rect 4552 7 4586 41
rect 4586 7 4598 41
rect 4546 -2 4598 7
rect 4610 41 4662 50
rect 4610 7 4624 41
rect 4624 7 4658 41
rect 4658 7 4662 41
rect 4610 -2 4662 7
rect 5666 75 5675 89
rect 5675 75 5709 89
rect 5709 75 5718 89
rect 5666 37 5718 75
rect 4253 -45 4262 -11
rect 4262 -45 4296 -11
rect 4296 -45 4305 -11
rect 4253 -46 4305 -45
rect 5265 -90 5317 -38
rect 4465 -120 4517 -111
rect 4465 -154 4471 -120
rect 4471 -154 4505 -120
rect 4505 -154 4517 -120
rect 4465 -163 4517 -154
rect 4529 -120 4581 -111
rect 4529 -154 4543 -120
rect 4543 -154 4577 -120
rect 4577 -154 4581 -120
rect 4529 -163 4581 -154
rect 4807 -119 4859 -110
rect 4871 -119 4923 -110
rect 4807 -153 4811 -119
rect 4811 -153 4859 -119
rect 4871 -153 4902 -119
rect 4902 -153 4923 -119
rect 4807 -162 4859 -153
rect 4871 -162 4923 -153
rect 5265 -154 5317 -102
rect 4363 -264 4415 -258
rect 4363 -298 4372 -264
rect 4372 -298 4406 -264
rect 4406 -298 4415 -264
rect 4363 -310 4415 -298
rect 4363 -339 4415 -322
rect 4363 -373 4372 -339
rect 4372 -373 4406 -339
rect 4406 -373 4415 -339
rect 5244 -264 5296 -212
rect 5244 -328 5296 -276
rect 4363 -374 4415 -373
rect 5666 -1 5675 25
rect 5675 -1 5709 25
rect 5709 -1 5718 25
rect 5666 -27 5718 -1
rect 3669 -794 3720 -760
rect 3720 -794 3721 -760
rect 3669 -796 3721 -794
rect 3601 -864 3653 -812
rect 3669 -864 3721 -812
rect 3601 -912 3604 -880
rect 3604 -912 3642 -880
rect 3642 -912 3653 -880
rect 3669 -912 3676 -880
rect 3676 -912 3714 -880
rect 3714 -912 3721 -880
rect 3601 -932 3653 -912
rect 3669 -932 3721 -912
<< metal2 >>
rect 3637 2365 3689 2371
rect 3885 2364 3937 2370
rect 3637 2312 3689 2313
tri 3689 2312 3706 2329 sw
rect 3386 2253 3392 2305
rect 3444 2253 3456 2305
rect 3508 2253 3514 2305
tri 3428 2249 3432 2253 ne
rect 3432 2249 3514 2253
tri 3432 2248 3433 2249 ne
rect 3433 2248 3514 2249
tri 3433 2219 3462 2248 ne
rect 703 2173 831 2179
rect 755 2121 831 2173
rect 703 2091 831 2121
rect 755 2039 831 2091
rect 703 2008 831 2039
rect 755 1956 831 2008
rect 703 1925 831 1956
rect 755 1873 831 1925
rect 125 1773 131 1825
rect 183 1773 195 1825
rect 247 1773 253 1825
rect 125 1725 253 1773
rect 125 1673 131 1725
rect 183 1673 195 1725
rect 247 1673 253 1725
rect 543 1774 549 1826
rect 601 1774 613 1826
rect 665 1774 671 1826
rect 543 385 671 1774
rect 703 1405 831 1873
rect 1713 2166 1841 2172
rect 1713 2114 1763 2166
rect 1815 2114 1841 2166
rect 1713 2084 1841 2114
rect 1713 2032 1763 2084
rect 1815 2032 1841 2084
rect 1713 2002 1841 2032
rect 1713 1950 1763 2002
rect 1815 1950 1841 2002
rect 1713 1919 1841 1950
rect 1713 1867 1763 1919
rect 1815 1867 1841 1919
rect 1036 1774 1042 1826
rect 1094 1774 1106 1826
rect 1158 1774 1164 1826
rect 1036 1565 1164 1774
rect 1036 1513 1042 1565
rect 1094 1513 1106 1565
rect 1158 1513 1164 1565
rect 1557 1773 1563 1825
rect 1615 1773 1627 1825
rect 1679 1773 1685 1825
rect 1557 1565 1685 1773
rect 1557 1513 1563 1565
rect 1615 1513 1627 1565
rect 1679 1513 1685 1565
rect 703 1353 709 1405
rect 761 1353 773 1405
rect 825 1353 831 1405
rect 703 945 831 1353
rect 1186 1433 1192 1485
rect 1244 1433 1256 1485
rect 1308 1433 1316 1485
tri 703 875 773 945 ne
rect 773 875 831 945
tri 831 875 955 999 sw
tri 773 848 800 875 ne
rect 800 848 955 875
tri 800 821 827 848 ne
rect 543 333 549 385
rect 601 333 613 385
rect 665 333 671 385
rect 543 289 671 333
rect 543 237 549 289
rect 601 237 613 289
rect 665 237 671 289
rect 827 70 955 848
rect 1186 289 1316 1433
rect 1713 1325 1841 1867
rect 1713 1273 1719 1325
rect 1771 1273 1783 1325
rect 1835 1273 1841 1325
rect 2075 2166 2127 2172
rect 2075 2084 2127 2114
rect 2075 2002 2127 2032
rect 2075 1919 2127 1950
rect 2075 1273 2127 1867
rect 2284 1773 2290 1825
rect 2342 1773 2354 1825
rect 2406 1773 2412 1825
rect 2284 1725 2412 1773
rect 2284 1673 2290 1725
rect 2342 1673 2354 1725
rect 2406 1673 2412 1725
rect 2500 1774 2506 1826
rect 2558 1774 2570 1826
rect 2622 1774 2628 1826
rect 2785 1774 2791 1826
rect 2843 1774 2855 1826
rect 2907 1774 2930 1826
rect 2500 1405 2628 1774
tri 2844 1740 2878 1774 ne
rect 2500 1353 2506 1405
rect 2558 1353 2570 1405
rect 2622 1353 2628 1405
rect 2722 1353 2728 1405
rect 2780 1353 2792 1405
rect 2844 1353 2850 1405
tri 2764 1325 2792 1353 ne
rect 2792 1325 2850 1353
tri 2127 1273 2133 1279 sw
rect 2588 1273 2594 1325
rect 2646 1273 2658 1325
rect 2710 1273 2716 1325
tri 2792 1319 2798 1325 ne
rect 2075 1245 2133 1273
tri 2133 1245 2161 1273 sw
rect 2075 1193 2081 1245
rect 2133 1193 2145 1245
rect 2197 1193 2203 1245
rect 1186 237 1192 289
rect 1244 237 1258 289
rect 1310 237 1316 289
rect 1869 333 1875 385
rect 1927 333 1939 385
rect 1991 333 1997 385
rect 1869 289 1997 333
rect 1869 237 1875 289
rect 1927 237 1939 289
rect 1991 237 1997 289
rect 879 18 903 70
rect 827 -19 955 18
rect 879 -71 903 -19
rect 827 -108 955 -71
rect 879 -160 903 -108
rect 827 -197 955 -160
rect 879 -249 903 -197
rect 827 -255 955 -249
rect -467 -638 -461 -586
rect -409 -638 -376 -586
rect -324 -638 -291 -586
rect -239 -638 -207 -586
rect -155 -638 -123 -586
rect -71 -638 1657 -586
rect -467 -696 1657 -638
rect -467 -748 -461 -696
rect -409 -748 -376 -696
rect -324 -748 -291 -696
rect -239 -748 -207 -696
rect -155 -748 -123 -696
rect -71 -748 1657 -696
rect 2588 -676 2716 1273
rect 2798 292 2850 1325
rect 2878 644 2930 1774
rect 2975 1774 2981 1826
rect 3033 1774 3045 1826
rect 3097 1774 3103 1826
rect 3230 1790 3236 1842
rect 3288 1790 3300 1842
rect 3352 1790 3358 1842
rect 2975 730 3027 1774
tri 3027 1740 3061 1774 nw
rect 3230 1759 3285 1790
tri 3285 1759 3316 1790 nw
rect 3230 848 3282 1759
tri 3282 1756 3285 1759 nw
tri 3459 1756 3462 1759 se
rect 3462 1756 3514 2248
rect 3637 2301 3706 2312
rect 3689 2300 3706 2301
tri 3706 2300 3718 2312 sw
rect 3885 2300 3937 2312
rect 3689 2295 3718 2300
tri 3718 2295 3723 2300 sw
rect 3689 2249 3749 2295
rect 3637 2248 3749 2249
tri 3749 2248 3796 2295 sw
rect 3637 2243 3796 2248
tri 3796 2243 3801 2248 sw
tri 3727 2231 3739 2243 ne
rect 3739 2231 3801 2243
tri 3801 2231 3813 2243 sw
tri 3739 2221 3749 2231 ne
rect 3749 2221 3813 2231
tri 3749 2209 3761 2221 ne
tri 3428 1725 3459 1756 se
rect 3459 1725 3514 1756
rect 3386 1673 3392 1725
rect 3444 1673 3456 1725
rect 3508 1673 3514 1725
rect 3601 2154 3721 2160
rect 3653 2102 3669 2154
rect 3601 2079 3721 2102
rect 3653 2027 3669 2079
rect 3601 2003 3721 2027
rect 3653 1951 3669 2003
tri 3282 848 3316 882 sw
rect 3230 796 3236 848
rect 3288 796 3300 848
rect 3352 796 3358 848
tri 3027 730 3061 764 sw
rect 2975 678 2981 730
rect 3033 678 3045 730
rect 3097 678 3103 730
rect 2878 580 2930 592
rect 2878 522 2930 528
tri 2850 292 2881 323 sw
rect 2798 291 2881 292
tri 2881 291 2882 292 sw
rect 2798 289 2882 291
tri 2882 289 2884 291 sw
rect 2798 237 2804 289
rect 2856 237 2868 289
rect 2920 237 2926 289
rect 3601 68 3721 1951
rect 3761 1193 3813 2221
rect 3885 1565 3937 2248
rect 4877 1673 4883 1725
rect 4935 1673 4947 1725
rect 4999 1673 5005 1725
tri 3937 1565 3971 1599 sw
rect 3885 1513 3891 1565
rect 3943 1513 3955 1565
rect 4007 1513 4013 1565
rect 4287 1433 4293 1485
rect 4345 1433 4357 1485
rect 4409 1433 4415 1485
tri 4329 1405 4357 1433 ne
rect 4357 1405 4415 1433
tri 4357 1399 4363 1405 ne
tri 3813 1193 3815 1195 sw
rect 3761 1161 3815 1193
tri 3815 1161 3847 1193 sw
rect 3761 1109 3767 1161
rect 3819 1109 3831 1161
rect 3883 1109 3889 1161
rect 3789 237 3795 289
rect 3847 237 3859 289
rect 3911 237 3979 289
rect 4177 237 4183 289
rect 4235 237 4247 289
rect 4299 237 4305 289
tri 3893 203 3927 237 ne
rect 3653 16 3669 68
rect 3601 1 3721 16
rect 3653 -51 3669 1
rect 3601 -66 3721 -51
rect 3927 70 3979 237
tri 4219 203 4253 237 ne
rect 3927 6 3979 18
rect 3927 -52 3979 -46
rect 4253 70 4305 237
rect 4253 6 4305 18
rect 4253 -52 4305 -46
rect 3653 -118 3669 -66
rect 3601 -133 3721 -118
rect 3653 -185 3669 -133
rect 3601 -200 3721 -185
rect 3653 -252 3669 -200
rect 3601 -268 3721 -252
rect 3653 -320 3669 -268
rect 3601 -336 3721 -320
rect 3653 -388 3669 -336
rect 4363 -258 4415 1405
rect 4570 1353 4576 1405
rect 4628 1353 4640 1405
rect 4692 1353 4698 1405
tri 4612 1319 4646 1353 ne
rect 4464 1193 4470 1245
rect 4522 1193 4534 1245
rect 4586 1193 4592 1245
tri 4506 1159 4540 1193 ne
rect 4459 547 4511 553
rect 4459 483 4511 495
rect 4459 -90 4511 431
rect 4540 50 4592 1193
rect 4646 292 4698 1353
tri 4698 292 4729 323 sw
rect 4646 291 4729 292
tri 4729 291 4730 292 sw
rect 4646 289 4730 291
tri 4730 289 4732 291 sw
rect 4646 237 4652 289
rect 4704 237 4716 289
rect 4768 237 4774 289
tri 4592 50 4629 87 sw
rect 4540 -2 4546 50
rect 4598 -2 4610 50
rect 4662 -2 4668 50
tri 4876 -77 4877 -76 se
rect 4877 -77 4929 1673
tri 4929 1639 4963 1673 nw
rect 5630 796 5636 848
rect 5688 796 5700 848
rect 5752 796 5758 848
tri 5672 762 5706 796 ne
rect 5474 678 5480 730
rect 5532 678 5544 730
rect 5596 678 5602 730
tri 5516 650 5544 678 ne
rect 5544 650 5602 678
rect 5371 598 5377 650
rect 5429 598 5441 650
rect 5493 598 5499 650
tri 5544 644 5550 650 ne
rect 5371 292 5499 598
rect 5189 239 5195 291
rect 5247 239 5259 291
rect 5311 239 5317 291
tri 5225 237 5227 239 ne
rect 5227 237 5317 239
tri 5227 199 5265 237 ne
tri 4511 -90 4524 -77 sw
tri 4863 -90 4876 -77 se
rect 4876 -90 4929 -77
rect 4459 -102 4524 -90
tri 4524 -102 4536 -90 sw
tri 4851 -102 4863 -90 se
rect 4863 -102 4929 -90
rect 4459 -110 4536 -102
tri 4536 -110 4544 -102 sw
tri 4843 -110 4851 -102 se
rect 4851 -110 4929 -102
rect 4459 -111 4544 -110
tri 4544 -111 4545 -110 sw
rect 4459 -163 4465 -111
rect 4517 -163 4529 -111
rect 4581 -163 4587 -111
rect 4801 -162 4807 -110
rect 4859 -162 4871 -110
rect 4923 -162 4929 -110
rect 5265 -38 5317 237
rect 5265 -102 5317 -90
rect 5265 -160 5317 -154
rect 5371 240 5377 292
rect 5429 240 5441 292
rect 5493 240 5499 292
rect 5550 289 5602 650
tri 5602 289 5636 323 sw
rect 5371 237 5454 240
tri 5454 237 5457 240 nw
rect 5550 237 5556 289
rect 5608 237 5620 289
rect 5672 237 5678 289
tri 5342 -206 5371 -177 se
rect 5371 -199 5423 237
tri 5423 206 5454 237 nw
tri 5684 153 5706 175 se
rect 5706 153 5758 796
tri 5666 135 5684 153 se
rect 5684 135 5718 153
rect 5666 89 5718 135
tri 5718 113 5758 153 nw
rect 5666 25 5718 37
rect 5666 -33 5718 -27
rect 5371 -206 5416 -199
tri 5416 -206 5423 -199 nw
rect 4363 -322 4415 -310
rect 5244 -212 5364 -206
rect 5296 -258 5364 -212
tri 5364 -258 5416 -206 nw
rect 5244 -276 5296 -264
tri 5296 -292 5330 -258 nw
rect 5244 -334 5296 -328
rect 4363 -380 4415 -374
rect 3601 -404 3721 -388
rect 3653 -456 3669 -404
rect 3601 -472 3721 -456
rect 3653 -524 3669 -472
rect 3601 -540 3721 -524
rect 3653 -592 3669 -540
rect 3601 -608 3721 -592
rect 3653 -660 3669 -608
tri 2716 -676 2720 -672 sw
rect 3601 -676 3721 -660
rect 2588 -706 2720 -676
tri 2720 -706 2750 -676 sw
rect 2588 -730 2758 -706
rect 2588 -782 2636 -730
rect 2688 -782 2700 -730
rect 2752 -782 2758 -730
rect 2588 -806 2758 -782
rect 3653 -728 3669 -676
rect 3601 -744 3721 -728
rect 3653 -796 3669 -744
rect 3601 -812 3721 -796
rect 3653 -864 3669 -812
rect 3601 -880 3721 -864
rect 3653 -932 3669 -880
rect 3601 -955 3721 -932
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1663361622
transform 1 0 3644 0 1 1921
box -46 24 399 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1663361622
transform -1 0 3826 0 1 1921
box 0 24 534 1116
use sky130_fd_pr__nfet_01v8__example_55959141808230  sky130_fd_pr__nfet_01v8__example_55959141808230_0
timestamp 1663361622
transform 1 0 4673 0 1 -802
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808230  sky130_fd_pr__nfet_01v8__example_55959141808230_1
timestamp 1663361622
transform 1 0 4985 0 1 -802
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808529  sky130_fd_pr__nfet_01v8__example_55959141808529_0
timestamp 1663361622
transform 1 0 4417 0 1 -802
box -1 0 201 1
use sky130_fd_pr__nfet_01v8__example_55959141808533  sky130_fd_pr__nfet_01v8__example_55959141808533_0
timestamp 1663361622
transform 1 0 5563 0 1 -802
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808533  sky130_fd_pr__nfet_01v8__example_55959141808533_1
timestamp 1663361622
transform 1 0 5407 0 1 -802
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808604  sky130_fd_pr__nfet_01v8__example_55959141808604_0
timestamp 1663361622
transform 1 0 3765 0 1 -802
box -1 0 161 1
use sky130_fd_pr__nfet_01v8__example_55959141808604  sky130_fd_pr__nfet_01v8__example_55959141808604_1
timestamp 1663361622
transform 1 0 4091 0 1 -802
box -1 0 161 1
use sky130_fd_pr__nfet_01v8__example_55959141808604  sky130_fd_pr__nfet_01v8__example_55959141808604_2
timestamp 1663361622
transform 1 0 1169 0 1 -802
box -1 0 161 1
use sky130_fd_pr__nfet_01v8__example_55959141808604  sky130_fd_pr__nfet_01v8__example_55959141808604_3
timestamp 1663361622
transform 1 0 3439 0 1 -802
box -1 0 161 1
use sky130_fd_pr__nfet_01v8__example_55959141808608  sky130_fd_pr__nfet_01v8__example_55959141808608_0
timestamp 1663361622
transform 1 0 4417 0 -1 213
box -1 0 809 1
use sky130_fd_pr__nfet_01v8__example_55959141808609  sky130_fd_pr__nfet_01v8__example_55959141808609_0
timestamp 1663361622
transform 1 0 2465 0 1 -802
box -1 0 809 1
use sky130_fd_pr__nfet_01v8__example_55959141808610  sky130_fd_pr__nfet_01v8__example_55959141808610_0
timestamp 1663361622
transform 1 0 1385 0 1 -802
box -1 0 1025 1
use sky130_fd_pr__nfet_01v8__example_55959141808610  sky130_fd_pr__nfet_01v8__example_55959141808610_1
timestamp 1663361622
transform 1 0 89 0 1 -802
box -1 0 1025 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_0
timestamp 1663361622
transform 1 0 1973 0 1 1865
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_1
timestamp 1663361622
transform 1 0 1661 0 1 1865
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_2
timestamp 1663361622
transform 1 0 119 0 1 1865
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_3
timestamp 1663361622
transform -1 0 1229 0 1 1865
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808548  sky130_fd_pr__pfet_01v8__example_55959141808548_0
timestamp 1663361622
transform 1 0 2817 0 1 1865
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808548  sky130_fd_pr__pfet_01v8__example_55959141808548_1
timestamp 1663361622
transform 1 0 2285 0 1 1865
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808548  sky130_fd_pr__pfet_01v8__example_55959141808548_2
timestamp 1663361622
transform 1 0 2973 0 1 1865
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808549  sky130_fd_pr__pfet_01v8__example_55959141808549_0
timestamp 1663361622
transform 1 0 2551 0 1 1865
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808611  sky130_fd_pr__pfet_01v8__example_55959141808611_0
timestamp 1663361622
transform 1 0 541 0 1 1865
box -1 0 161 1
use sky130_fd_pr__pfet_01v8__example_55959141808611  sky130_fd_pr__pfet_01v8__example_55959141808611_1
timestamp 1663361622
transform -1 0 1605 0 1 1865
box -1 0 161 1
use sky130_fd_pr__pfet_01v8__example_55959141808611  sky130_fd_pr__pfet_01v8__example_55959141808611_2
timestamp 1663361622
transform 1 0 757 0 1 1865
box -1 0 161 1
<< labels >>
flabel metal2 s 5717 586 5750 748 3 FreeSans 200 0 0 0 OUT
port 1 nsew
flabel metal2 s 5553 502 5593 628 3 FreeSans 200 0 0 0 OUT_N
port 2 nsew
flabel metal1 s 885 1677 973 1720 3 FreeSans 200 0 0 0 MODE_NORMAL_N
port 3 nsew
flabel metal1 s 284 350 354 381 3 FreeSans 200 0 0 0 IN_H
port 4 nsew
flabel metal1 s 272 1442 346 1478 3 FreeSans 200 0 0 0 IN_VT
port 5 nsew
flabel metal1 s 3646 2270 3677 2350 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 6 nsew
flabel metal1 s 4476 -152 4570 -123 3 FreeSans 200 0 0 0 VTRIP_SEL_H_N
port 7 nsew
flabel metal1 s 96 2865 297 3006 3 FreeSans 200 0 0 0 VDDIO_Q
port 8 nsew
flabel metal1 s 84 -1123 481 -913 3 FreeSans 200 0 0 0 VSSD
port 9 nsew
flabel comment s 400 1545 400 1545 0 FreeSans 200 0 0 0 MODE_NORMAL_CMOS_H_N
flabel comment s 625 1704 625 1704 0 FreeSans 200 0 0 0 MODE_NORMAL_N
flabel comment s 2754 1708 2754 1708 0 FreeSans 200 0 0 0 MODE_NORMAL_N
flabel comment s 400 1462 400 1462 0 FreeSans 200 0 0 0 IN_VT
<< properties >>
string GDS_END 45533758
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 45411946
<< end >>
