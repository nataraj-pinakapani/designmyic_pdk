/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/cdl/sky130_fd_io/sky130_ef_io.cdl