/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/lef/sky130_fd_sc_hd/sky130_ef_sc_hd.lef