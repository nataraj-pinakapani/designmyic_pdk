magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1907 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 423 47 453 177
rect 507 47 537 177
rect 591 47 621 177
rect 775 47 805 177
rect 859 47 889 177
rect 943 47 973 177
rect 1027 47 1057 177
rect 1111 47 1141 177
rect 1211 47 1241 177
rect 1295 47 1325 177
rect 1379 47 1409 177
rect 1463 47 1493 177
rect 1547 47 1577 177
rect 1631 47 1661 177
rect 1715 47 1745 177
rect 1799 47 1829 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 523 297 553 497
rect 607 297 637 497
rect 691 297 721 497
rect 775 297 805 497
rect 859 297 889 497
rect 943 297 973 497
rect 1027 297 1057 497
rect 1111 297 1141 497
rect 1211 297 1241 497
rect 1295 297 1325 497
rect 1379 297 1409 497
rect 1463 297 1493 497
rect 1547 297 1577 497
rect 1631 297 1661 497
rect 1715 297 1745 497
rect 1799 297 1829 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 423 177
rect 365 61 375 95
rect 409 61 423 95
rect 365 47 423 61
rect 453 95 507 177
rect 453 61 463 95
rect 497 61 507 95
rect 453 47 507 61
rect 537 169 591 177
rect 537 135 547 169
rect 581 135 591 169
rect 537 47 591 135
rect 621 95 775 177
rect 621 61 631 95
rect 665 61 731 95
rect 765 61 775 95
rect 621 47 775 61
rect 805 163 859 177
rect 805 129 815 163
rect 849 129 859 163
rect 805 47 859 129
rect 889 95 943 177
rect 889 61 899 95
rect 933 61 943 95
rect 889 47 943 61
rect 973 163 1027 177
rect 973 129 983 163
rect 1017 129 1027 163
rect 973 47 1027 129
rect 1057 95 1111 177
rect 1057 61 1067 95
rect 1101 61 1111 95
rect 1057 47 1111 61
rect 1141 95 1211 177
rect 1141 61 1167 95
rect 1201 61 1211 95
rect 1141 47 1211 61
rect 1241 95 1295 177
rect 1241 61 1251 95
rect 1285 61 1295 95
rect 1241 47 1295 61
rect 1325 163 1379 177
rect 1325 129 1335 163
rect 1369 129 1379 163
rect 1325 47 1379 129
rect 1409 95 1463 177
rect 1409 61 1419 95
rect 1453 61 1463 95
rect 1409 47 1463 61
rect 1493 163 1547 177
rect 1493 129 1503 163
rect 1537 129 1547 163
rect 1493 47 1547 129
rect 1577 163 1631 177
rect 1577 129 1587 163
rect 1621 129 1631 163
rect 1577 95 1631 129
rect 1577 61 1587 95
rect 1621 61 1631 95
rect 1577 47 1631 61
rect 1661 95 1715 177
rect 1661 61 1671 95
rect 1705 61 1715 95
rect 1661 47 1715 61
rect 1745 163 1799 177
rect 1745 129 1755 163
rect 1789 129 1799 163
rect 1745 95 1799 129
rect 1745 61 1755 95
rect 1789 61 1799 95
rect 1745 47 1799 61
rect 1829 163 1881 177
rect 1829 129 1839 163
rect 1873 129 1881 163
rect 1829 95 1881 129
rect 1829 61 1839 95
rect 1873 61 1881 95
rect 1829 47 1881 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 409 167 497
rect 113 375 123 409
rect 157 375 167 409
rect 113 341 167 375
rect 113 307 123 341
rect 157 307 167 341
rect 113 297 167 307
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 297 251 375
rect 281 409 335 497
rect 281 375 291 409
rect 325 375 335 409
rect 281 341 335 375
rect 281 307 291 341
rect 325 307 335 341
rect 281 297 335 307
rect 365 479 417 497
rect 365 445 375 479
rect 409 445 417 479
rect 365 411 417 445
rect 365 377 375 411
rect 409 377 417 411
rect 365 343 417 377
rect 365 309 375 343
rect 409 309 417 343
rect 365 297 417 309
rect 471 477 523 497
rect 471 443 479 477
rect 513 443 523 477
rect 471 409 523 443
rect 471 375 479 409
rect 513 375 523 409
rect 471 297 523 375
rect 553 409 607 497
rect 553 375 563 409
rect 597 375 607 409
rect 553 341 607 375
rect 553 307 563 341
rect 597 307 607 341
rect 553 297 607 307
rect 637 477 691 497
rect 637 443 647 477
rect 681 443 691 477
rect 637 297 691 443
rect 721 409 775 497
rect 721 375 731 409
rect 765 375 775 409
rect 721 297 775 375
rect 805 477 859 497
rect 805 443 815 477
rect 849 443 859 477
rect 805 297 859 443
rect 889 409 943 497
rect 889 375 899 409
rect 933 375 943 409
rect 889 297 943 375
rect 973 477 1027 497
rect 973 443 983 477
rect 1017 443 1027 477
rect 973 297 1027 443
rect 1057 409 1111 497
rect 1057 375 1067 409
rect 1101 375 1111 409
rect 1057 297 1111 375
rect 1141 477 1211 497
rect 1141 443 1159 477
rect 1193 443 1211 477
rect 1141 409 1211 443
rect 1141 375 1159 409
rect 1193 375 1211 409
rect 1141 297 1211 375
rect 1241 477 1295 497
rect 1241 443 1251 477
rect 1285 443 1295 477
rect 1241 297 1295 443
rect 1325 409 1379 497
rect 1325 375 1335 409
rect 1369 375 1379 409
rect 1325 297 1379 375
rect 1409 477 1463 497
rect 1409 443 1419 477
rect 1453 443 1463 477
rect 1409 297 1463 443
rect 1493 409 1547 497
rect 1493 375 1503 409
rect 1537 375 1547 409
rect 1493 297 1547 375
rect 1577 477 1631 497
rect 1577 443 1587 477
rect 1621 443 1631 477
rect 1577 297 1631 443
rect 1661 477 1715 497
rect 1661 443 1671 477
rect 1705 443 1715 477
rect 1661 409 1715 443
rect 1661 375 1671 409
rect 1705 375 1715 409
rect 1661 297 1715 375
rect 1745 477 1799 497
rect 1745 443 1755 477
rect 1789 443 1799 477
rect 1745 409 1799 443
rect 1745 375 1755 409
rect 1789 375 1799 409
rect 1745 297 1799 375
rect 1829 477 1888 497
rect 1829 443 1839 477
rect 1873 443 1888 477
rect 1829 409 1888 443
rect 1829 375 1839 409
rect 1873 375 1888 409
rect 1829 341 1888 375
rect 1829 307 1839 341
rect 1873 307 1888 341
rect 1829 297 1888 307
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 463 61 497 95
rect 547 135 581 169
rect 631 61 665 95
rect 731 61 765 95
rect 815 129 849 163
rect 899 61 933 95
rect 983 129 1017 163
rect 1067 61 1101 95
rect 1167 61 1201 95
rect 1251 61 1285 95
rect 1335 129 1369 163
rect 1419 61 1453 95
rect 1503 129 1537 163
rect 1587 129 1621 163
rect 1587 61 1621 95
rect 1671 61 1705 95
rect 1755 129 1789 163
rect 1755 61 1789 95
rect 1839 129 1873 163
rect 1839 61 1873 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 375 157 409
rect 123 307 157 341
rect 207 443 241 477
rect 207 375 241 409
rect 291 375 325 409
rect 291 307 325 341
rect 375 445 409 479
rect 375 377 409 411
rect 375 309 409 343
rect 479 443 513 477
rect 479 375 513 409
rect 563 375 597 409
rect 563 307 597 341
rect 647 443 681 477
rect 731 375 765 409
rect 815 443 849 477
rect 899 375 933 409
rect 983 443 1017 477
rect 1067 375 1101 409
rect 1159 443 1193 477
rect 1159 375 1193 409
rect 1251 443 1285 477
rect 1335 375 1369 409
rect 1419 443 1453 477
rect 1503 375 1537 409
rect 1587 443 1621 477
rect 1671 443 1705 477
rect 1671 375 1705 409
rect 1755 443 1789 477
rect 1755 375 1789 409
rect 1839 443 1873 477
rect 1839 375 1873 409
rect 1839 307 1873 341
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 523 497 553 523
rect 607 497 637 523
rect 691 497 721 523
rect 775 497 805 523
rect 859 497 889 523
rect 943 497 973 523
rect 1027 497 1057 523
rect 1111 497 1141 523
rect 1211 497 1241 523
rect 1295 497 1325 523
rect 1379 497 1409 523
rect 1463 497 1493 523
rect 1547 497 1577 523
rect 1631 497 1661 523
rect 1715 497 1745 523
rect 1799 497 1829 523
rect 83 265 113 297
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 523 265 553 297
rect 607 265 637 297
rect 691 265 721 297
rect 775 265 805 297
rect 859 265 889 297
rect 943 265 973 297
rect 1027 265 1057 297
rect 1111 265 1141 297
rect 1211 265 1241 297
rect 1295 265 1325 297
rect 1379 265 1409 297
rect 1463 265 1493 297
rect 1547 265 1577 297
rect 65 249 365 265
rect 65 215 81 249
rect 115 215 149 249
rect 183 215 217 249
rect 251 215 365 249
rect 65 199 365 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 423 249 727 265
rect 423 215 683 249
rect 717 215 727 249
rect 423 199 727 215
rect 775 249 1057 265
rect 775 215 803 249
rect 837 215 871 249
rect 905 215 939 249
rect 973 215 1007 249
rect 1041 215 1057 249
rect 775 199 1057 215
rect 1099 249 1153 265
rect 1099 215 1109 249
rect 1143 215 1153 249
rect 1099 199 1153 215
rect 1199 249 1253 265
rect 1199 215 1209 249
rect 1243 215 1253 249
rect 1199 199 1253 215
rect 1295 249 1577 265
rect 1295 215 1311 249
rect 1345 215 1379 249
rect 1413 215 1447 249
rect 1481 215 1515 249
rect 1549 215 1577 249
rect 1295 199 1577 215
rect 423 177 453 199
rect 507 177 537 199
rect 591 177 621 199
rect 775 177 805 199
rect 859 177 889 199
rect 943 177 973 199
rect 1027 177 1057 199
rect 1111 177 1141 199
rect 1211 177 1241 199
rect 1295 177 1325 199
rect 1379 177 1409 199
rect 1463 177 1493 199
rect 1547 177 1577 199
rect 1631 265 1661 297
rect 1715 265 1745 297
rect 1799 265 1829 297
rect 1631 249 1838 265
rect 1631 215 1647 249
rect 1681 215 1715 249
rect 1749 215 1783 249
rect 1817 215 1838 249
rect 1631 199 1838 215
rect 1631 177 1661 199
rect 1715 177 1745 199
rect 1799 177 1829 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 423 21 453 47
rect 507 21 537 47
rect 591 21 621 47
rect 775 21 805 47
rect 859 21 889 47
rect 943 21 973 47
rect 1027 21 1057 47
rect 1111 21 1141 47
rect 1211 21 1241 47
rect 1295 21 1325 47
rect 1379 21 1409 47
rect 1463 21 1493 47
rect 1547 21 1577 47
rect 1631 21 1661 47
rect 1715 21 1745 47
rect 1799 21 1829 47
<< polycont >>
rect 81 215 115 249
rect 149 215 183 249
rect 217 215 251 249
rect 683 215 717 249
rect 803 215 837 249
rect 871 215 905 249
rect 939 215 973 249
rect 1007 215 1041 249
rect 1109 215 1143 249
rect 1209 215 1243 249
rect 1311 215 1345 249
rect 1379 215 1413 249
rect 1447 215 1481 249
rect 1515 215 1549 249
rect 1647 215 1681 249
rect 1715 215 1749 249
rect 1783 215 1817 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 18 479 425 493
rect 18 477 375 479
rect 18 443 39 477
rect 73 459 207 477
rect 73 443 81 459
rect 18 409 81 443
rect 199 443 207 459
rect 241 459 375 477
rect 241 443 249 459
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 18 307 39 341
rect 73 307 81 341
rect 18 289 81 307
rect 115 409 165 425
rect 115 375 123 409
rect 157 375 165 409
rect 115 341 165 375
rect 199 409 249 443
rect 409 445 425 479
rect 199 375 207 409
rect 241 375 249 409
rect 199 357 249 375
rect 283 409 333 425
rect 283 375 291 409
rect 325 375 333 409
rect 115 307 123 341
rect 157 323 165 341
rect 283 341 333 375
rect 283 323 291 341
rect 157 307 291 323
rect 325 323 333 341
rect 375 411 425 445
rect 409 377 425 411
rect 375 343 425 377
rect 463 477 1201 493
rect 463 443 479 477
rect 513 443 647 477
rect 681 443 815 477
rect 849 443 983 477
rect 1017 443 1159 477
rect 1193 443 1201 477
rect 1235 477 1637 527
rect 1235 443 1251 477
rect 1285 443 1419 477
rect 1453 443 1587 477
rect 1621 443 1637 477
rect 1671 477 1705 493
rect 463 409 513 443
rect 1151 409 1201 443
rect 1671 409 1705 443
rect 1755 477 1789 527
rect 1755 409 1789 443
rect 463 375 479 409
rect 463 359 513 375
rect 547 375 563 409
rect 597 375 731 409
rect 765 375 899 409
rect 933 375 1067 409
rect 1101 375 1117 409
rect 547 367 1117 375
rect 1151 375 1159 409
rect 1193 375 1335 409
rect 1369 375 1503 409
rect 1537 375 1671 409
rect 1705 375 1721 409
rect 325 307 341 323
rect 115 289 341 307
rect 409 323 425 343
rect 547 341 606 367
rect 1151 357 1721 375
rect 1755 359 1789 375
rect 1831 477 1881 493
rect 1831 443 1839 477
rect 1873 443 1881 477
rect 1831 409 1881 443
rect 1831 375 1839 409
rect 1873 375 1881 409
rect 547 323 563 341
rect 409 309 563 323
rect 375 307 563 309
rect 597 307 606 341
rect 1687 323 1721 357
rect 1831 341 1881 375
rect 1831 323 1839 341
rect 375 289 606 307
rect 719 289 1159 323
rect 301 255 341 289
rect 719 265 753 289
rect 18 249 267 255
rect 18 215 81 249
rect 115 215 149 249
rect 183 215 217 249
rect 251 215 267 249
rect 301 219 649 255
rect 301 181 341 219
rect 23 163 73 179
rect 23 129 39 163
rect 23 95 73 129
rect 23 61 39 95
rect 23 17 73 61
rect 107 163 341 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 129 341 163
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 169 581 185
rect 375 135 547 169
rect 375 129 581 135
rect 615 164 649 219
rect 683 249 753 265
rect 717 215 753 249
rect 683 199 753 215
rect 787 249 1057 255
rect 787 215 803 249
rect 837 215 871 249
rect 905 215 939 249
rect 973 215 1007 249
rect 1041 215 1057 249
rect 1093 249 1159 289
rect 1093 215 1109 249
rect 1143 215 1159 249
rect 1193 289 1653 323
rect 1687 307 1839 323
rect 1873 307 1881 341
rect 1687 289 1881 307
rect 1193 249 1259 289
rect 1619 255 1653 289
rect 1193 215 1209 249
rect 1243 215 1259 249
rect 1295 249 1577 255
rect 1295 215 1311 249
rect 1345 215 1379 249
rect 1413 215 1447 249
rect 1481 215 1515 249
rect 1549 215 1577 249
rect 1619 249 1915 255
rect 1619 215 1647 249
rect 1681 215 1715 249
rect 1749 215 1783 249
rect 1817 215 1915 249
rect 787 199 1057 215
rect 1102 164 1292 181
rect 615 163 1553 164
rect 615 129 815 163
rect 849 129 983 163
rect 1017 147 1335 163
rect 1017 129 1136 147
rect 1258 129 1335 147
rect 1369 129 1503 163
rect 1537 129 1553 163
rect 1587 163 1805 181
rect 1621 145 1755 163
rect 1621 129 1637 145
rect 375 95 409 129
rect 547 119 581 129
rect 1167 95 1201 111
rect 1587 95 1637 129
rect 1739 129 1755 145
rect 1789 129 1805 163
rect 375 17 409 61
rect 447 61 463 95
rect 497 85 522 95
rect 607 85 631 95
rect 497 61 631 85
rect 665 61 731 95
rect 765 61 899 95
rect 933 61 1067 95
rect 1101 61 1117 95
rect 447 51 1117 61
rect 1167 17 1201 61
rect 1235 61 1251 95
rect 1285 61 1419 95
rect 1453 61 1587 95
rect 1621 61 1637 95
rect 1235 51 1637 61
rect 1671 95 1705 111
rect 1671 17 1705 61
rect 1739 95 1805 129
rect 1739 61 1755 95
rect 1789 61 1805 95
rect 1739 51 1805 61
rect 1839 163 1873 181
rect 1839 95 1873 129
rect 1839 17 1873 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 1690 221 1724 255 0 FreeSans 400 180 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 400 180 0 0 Y
port 10 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel locali s 1414 221 1448 255 0 FreeSans 400 180 0 0 A1
port 1 nsew signal input
flabel locali s 770 289 804 323 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 a221oi_4
rlabel metal1 s 0 -48 1932 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 3687728
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 3674506
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 48.300 0.000 
<< end >>
