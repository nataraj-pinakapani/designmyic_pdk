magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 5702 9167 6448 12639
rect 5839 9166 6373 9167
<< pwell >>
rect -10296 8021 -9842 8027
rect -10296 7936 -9590 8021
rect -10542 7378 -9590 7936
rect -10296 7375 -9590 7378
rect -9726 7182 -9590 7375
rect -10492 7007 -9590 7182
rect -10492 6824 -9816 7007
rect -10492 6670 -1845 6824
rect -10492 6644 -5512 6670
rect -10638 6392 -5512 6644
rect -10373 5938 -10095 6190
<< mvnmos >>
rect -10516 7457 -10432 7857
rect -10217 7401 -10097 8001
rect -10041 7401 -9921 8001
rect -9700 7542 -9616 7942
rect -9700 7086 -9616 7486
rect -10559 6418 -9759 6618
rect -9703 6418 -8103 6618
rect -8047 6418 -6447 6618
rect -6391 6418 -5591 6618
rect -10294 5964 -10174 6164
<< mvpmos >>
rect 5821 12433 5941 12573
rect 6179 12433 6299 12573
rect 5782 12059 6382 12179
rect 5782 11883 6382 12003
rect 5782 11707 6382 11827
rect 5782 11451 6382 11651
rect 5782 11195 6382 11395
rect 5782 10939 6382 11139
rect 5782 10683 6382 10883
rect 5782 10427 6382 10627
rect 5782 10171 6382 10371
rect 5782 9915 6382 10115
rect 5782 9659 6382 9859
rect 5958 9232 6078 9432
rect 6134 9232 6254 9432
<< mvndiff >>
rect -10270 7989 -10217 8001
rect -10270 7955 -10262 7989
rect -10228 7955 -10217 7989
rect -10270 7921 -10217 7955
rect -10516 7902 -10432 7910
rect -10516 7868 -10478 7902
rect -10444 7868 -10432 7902
rect -10516 7857 -10432 7868
rect -10270 7887 -10262 7921
rect -10228 7887 -10217 7921
rect -10270 7853 -10217 7887
rect -10270 7819 -10262 7853
rect -10228 7819 -10217 7853
rect -10270 7785 -10217 7819
rect -10270 7751 -10262 7785
rect -10228 7751 -10217 7785
rect -10270 7717 -10217 7751
rect -10270 7683 -10262 7717
rect -10228 7683 -10217 7717
rect -10270 7649 -10217 7683
rect -10270 7615 -10262 7649
rect -10228 7615 -10217 7649
rect -10270 7581 -10217 7615
rect -10270 7547 -10262 7581
rect -10228 7547 -10217 7581
rect -10270 7513 -10217 7547
rect -10270 7479 -10262 7513
rect -10228 7479 -10217 7513
rect -10516 7446 -10432 7457
rect -10516 7412 -10478 7446
rect -10444 7412 -10432 7446
rect -10516 7404 -10432 7412
rect -10270 7401 -10217 7479
rect -10097 7989 -10041 8001
rect -10097 7955 -10086 7989
rect -10052 7955 -10041 7989
rect -10097 7921 -10041 7955
rect -10097 7887 -10086 7921
rect -10052 7887 -10041 7921
rect -10097 7853 -10041 7887
rect -10097 7819 -10086 7853
rect -10052 7819 -10041 7853
rect -10097 7785 -10041 7819
rect -10097 7751 -10086 7785
rect -10052 7751 -10041 7785
rect -10097 7717 -10041 7751
rect -10097 7683 -10086 7717
rect -10052 7683 -10041 7717
rect -10097 7649 -10041 7683
rect -10097 7615 -10086 7649
rect -10052 7615 -10041 7649
rect -10097 7581 -10041 7615
rect -10097 7547 -10086 7581
rect -10052 7547 -10041 7581
rect -10097 7513 -10041 7547
rect -10097 7479 -10086 7513
rect -10052 7479 -10041 7513
rect -10097 7401 -10041 7479
rect -9921 7989 -9868 8001
rect -9921 7955 -9910 7989
rect -9876 7955 -9868 7989
rect -9921 7921 -9868 7955
rect -9700 7987 -9616 7995
rect -9700 7953 -9662 7987
rect -9628 7953 -9616 7987
rect -9700 7942 -9616 7953
rect -9921 7887 -9910 7921
rect -9876 7887 -9868 7921
rect -9921 7853 -9868 7887
rect -9921 7819 -9910 7853
rect -9876 7819 -9868 7853
rect -9921 7785 -9868 7819
rect -9921 7751 -9910 7785
rect -9876 7751 -9868 7785
rect -9921 7717 -9868 7751
rect -9921 7683 -9910 7717
rect -9876 7683 -9868 7717
rect -9921 7649 -9868 7683
rect -9921 7615 -9910 7649
rect -9876 7615 -9868 7649
rect -9921 7581 -9868 7615
rect -9921 7547 -9910 7581
rect -9876 7547 -9868 7581
rect -9921 7513 -9868 7547
rect -9921 7479 -9910 7513
rect -9876 7479 -9868 7513
rect -9700 7531 -9616 7542
rect -9700 7497 -9662 7531
rect -9628 7497 -9616 7531
rect -9700 7486 -9616 7497
rect -9921 7401 -9868 7479
rect -9700 7075 -9616 7086
rect -9700 7041 -9662 7075
rect -9628 7041 -9616 7075
rect -9700 7033 -9616 7041
rect -10612 6606 -10559 6618
rect -10612 6572 -10604 6606
rect -10570 6572 -10559 6606
rect -10612 6538 -10559 6572
rect -10612 6504 -10604 6538
rect -10570 6504 -10559 6538
rect -10612 6470 -10559 6504
rect -10612 6436 -10604 6470
rect -10570 6436 -10559 6470
rect -10612 6418 -10559 6436
rect -9759 6606 -9703 6618
rect -9759 6572 -9748 6606
rect -9714 6572 -9703 6606
rect -9759 6538 -9703 6572
rect -9759 6504 -9748 6538
rect -9714 6504 -9703 6538
rect -9759 6470 -9703 6504
rect -9759 6436 -9748 6470
rect -9714 6436 -9703 6470
rect -9759 6418 -9703 6436
rect -8103 6606 -8047 6618
rect -8103 6572 -8092 6606
rect -8058 6572 -8047 6606
rect -8103 6538 -8047 6572
rect -8103 6504 -8092 6538
rect -8058 6504 -8047 6538
rect -8103 6470 -8047 6504
rect -8103 6436 -8092 6470
rect -8058 6436 -8047 6470
rect -8103 6418 -8047 6436
rect -6447 6606 -6391 6618
rect -6447 6572 -6436 6606
rect -6402 6572 -6391 6606
rect -6447 6538 -6391 6572
rect -6447 6504 -6436 6538
rect -6402 6504 -6391 6538
rect -6447 6470 -6391 6504
rect -6447 6436 -6436 6470
rect -6402 6436 -6391 6470
rect -6447 6418 -6391 6436
rect -5591 6606 -5538 6618
rect -5591 6572 -5580 6606
rect -5546 6572 -5538 6606
rect -5591 6538 -5538 6572
rect -5591 6504 -5580 6538
rect -5546 6504 -5538 6538
rect -5591 6470 -5538 6504
rect -5591 6436 -5580 6470
rect -5546 6436 -5538 6470
rect -5591 6418 -5538 6436
rect -10347 6146 -10294 6164
rect -10347 6112 -10339 6146
rect -10305 6112 -10294 6146
rect -10347 6078 -10294 6112
rect -10347 6044 -10339 6078
rect -10305 6044 -10294 6078
rect -10347 6010 -10294 6044
rect -10347 5976 -10339 6010
rect -10305 5976 -10294 6010
rect -10347 5964 -10294 5976
rect -10174 6146 -10121 6164
rect -10174 6112 -10163 6146
rect -10129 6112 -10121 6146
rect -10174 6078 -10121 6112
rect -10174 6044 -10163 6078
rect -10129 6044 -10121 6078
rect -10174 6010 -10121 6044
rect -10174 5976 -10163 6010
rect -10129 5976 -10121 6010
rect -10174 5964 -10121 5976
<< mvpdiff >>
rect 5768 12547 5821 12573
rect 5768 12513 5776 12547
rect 5810 12513 5821 12547
rect 5768 12479 5821 12513
rect 5768 12445 5776 12479
rect 5810 12445 5821 12479
rect 5768 12433 5821 12445
rect 5941 12547 5994 12573
rect 5941 12513 5952 12547
rect 5986 12513 5994 12547
rect 5941 12479 5994 12513
rect 5941 12445 5952 12479
rect 5986 12445 5994 12479
rect 5941 12433 5994 12445
rect 6126 12547 6179 12573
rect 6126 12513 6134 12547
rect 6168 12513 6179 12547
rect 6126 12479 6179 12513
rect 6126 12445 6134 12479
rect 6168 12445 6179 12479
rect 6126 12433 6179 12445
rect 6299 12547 6352 12573
rect 6299 12513 6310 12547
rect 6344 12513 6352 12547
rect 6299 12479 6352 12513
rect 6299 12445 6310 12479
rect 6344 12445 6352 12479
rect 6299 12433 6352 12445
rect 5782 12224 6382 12232
rect 5782 12190 5860 12224
rect 5894 12190 5928 12224
rect 5962 12190 5996 12224
rect 6030 12190 6064 12224
rect 6098 12190 6132 12224
rect 6166 12190 6200 12224
rect 6234 12190 6268 12224
rect 6302 12190 6336 12224
rect 6370 12190 6382 12224
rect 5782 12179 6382 12190
rect 5782 12048 6382 12059
rect 5782 12014 5860 12048
rect 5894 12014 5928 12048
rect 5962 12014 5996 12048
rect 6030 12014 6064 12048
rect 6098 12014 6132 12048
rect 6166 12014 6200 12048
rect 6234 12014 6268 12048
rect 6302 12014 6336 12048
rect 6370 12014 6382 12048
rect 5782 12003 6382 12014
rect 5782 11872 6382 11883
rect 5782 11838 5860 11872
rect 5894 11838 5928 11872
rect 5962 11838 5996 11872
rect 6030 11838 6064 11872
rect 6098 11838 6132 11872
rect 6166 11838 6200 11872
rect 6234 11838 6268 11872
rect 6302 11838 6336 11872
rect 6370 11838 6382 11872
rect 5782 11827 6382 11838
rect 5782 11696 6382 11707
rect 5782 11662 5860 11696
rect 5894 11662 5928 11696
rect 5962 11662 5996 11696
rect 6030 11662 6064 11696
rect 6098 11662 6132 11696
rect 6166 11662 6200 11696
rect 6234 11662 6268 11696
rect 6302 11662 6336 11696
rect 6370 11662 6382 11696
rect 5782 11651 6382 11662
rect 5782 11440 6382 11451
rect 5782 11406 5860 11440
rect 5894 11406 5928 11440
rect 5962 11406 5996 11440
rect 6030 11406 6064 11440
rect 6098 11406 6132 11440
rect 6166 11406 6200 11440
rect 6234 11406 6268 11440
rect 6302 11406 6336 11440
rect 6370 11406 6382 11440
rect 5782 11395 6382 11406
rect 5782 11184 6382 11195
rect 5782 11150 5860 11184
rect 5894 11150 5928 11184
rect 5962 11150 5996 11184
rect 6030 11150 6064 11184
rect 6098 11150 6132 11184
rect 6166 11150 6200 11184
rect 6234 11150 6268 11184
rect 6302 11150 6336 11184
rect 6370 11150 6382 11184
rect 5782 11139 6382 11150
rect 5782 10928 6382 10939
rect 5782 10894 5860 10928
rect 5894 10894 5928 10928
rect 5962 10894 5996 10928
rect 6030 10894 6064 10928
rect 6098 10894 6132 10928
rect 6166 10894 6200 10928
rect 6234 10894 6268 10928
rect 6302 10894 6336 10928
rect 6370 10894 6382 10928
rect 5782 10883 6382 10894
rect 5782 10672 6382 10683
rect 5782 10638 5860 10672
rect 5894 10638 5928 10672
rect 5962 10638 5996 10672
rect 6030 10638 6064 10672
rect 6098 10638 6132 10672
rect 6166 10638 6200 10672
rect 6234 10638 6268 10672
rect 6302 10638 6336 10672
rect 6370 10638 6382 10672
rect 5782 10627 6382 10638
rect 5782 10416 6382 10427
rect 5782 10382 5860 10416
rect 5894 10382 5928 10416
rect 5962 10382 5996 10416
rect 6030 10382 6064 10416
rect 6098 10382 6132 10416
rect 6166 10382 6200 10416
rect 6234 10382 6268 10416
rect 6302 10382 6336 10416
rect 6370 10382 6382 10416
rect 5782 10371 6382 10382
rect 5782 10160 6382 10171
rect 5782 10126 5860 10160
rect 5894 10126 5928 10160
rect 5962 10126 5996 10160
rect 6030 10126 6064 10160
rect 6098 10126 6132 10160
rect 6166 10126 6200 10160
rect 6234 10126 6268 10160
rect 6302 10126 6336 10160
rect 6370 10126 6382 10160
rect 5782 10115 6382 10126
rect 5782 9904 6382 9915
rect 5782 9870 5860 9904
rect 5894 9870 5928 9904
rect 5962 9870 5996 9904
rect 6030 9870 6064 9904
rect 6098 9870 6132 9904
rect 6166 9870 6200 9904
rect 6234 9870 6268 9904
rect 6302 9870 6336 9904
rect 6370 9870 6382 9904
rect 5782 9859 6382 9870
rect 5782 9648 6382 9659
rect 5782 9614 5860 9648
rect 5894 9614 5928 9648
rect 5962 9614 5996 9648
rect 6030 9614 6064 9648
rect 6098 9614 6132 9648
rect 6166 9614 6200 9648
rect 6234 9614 6268 9648
rect 6302 9614 6336 9648
rect 6370 9614 6382 9648
rect 5782 9606 6382 9614
rect 5905 9420 5958 9432
rect 5905 9386 5913 9420
rect 5947 9386 5958 9420
rect 5905 9352 5958 9386
rect 5905 9318 5913 9352
rect 5947 9318 5958 9352
rect 5905 9284 5958 9318
rect 5905 9250 5913 9284
rect 5947 9250 5958 9284
rect 5905 9232 5958 9250
rect 6078 9420 6134 9432
rect 6078 9386 6089 9420
rect 6123 9386 6134 9420
rect 6078 9352 6134 9386
rect 6078 9318 6089 9352
rect 6123 9318 6134 9352
rect 6078 9284 6134 9318
rect 6078 9250 6089 9284
rect 6123 9250 6134 9284
rect 6078 9232 6134 9250
rect 6254 9420 6307 9432
rect 6254 9386 6265 9420
rect 6299 9386 6307 9420
rect 6254 9352 6307 9386
rect 6254 9318 6265 9352
rect 6299 9318 6307 9352
rect 6254 9284 6307 9318
rect 6254 9250 6265 9284
rect 6299 9250 6307 9284
rect 6254 9232 6307 9250
<< mvndiffc >>
rect -10262 7955 -10228 7989
rect -10478 7868 -10444 7902
rect -10262 7887 -10228 7921
rect -10262 7819 -10228 7853
rect -10262 7751 -10228 7785
rect -10262 7683 -10228 7717
rect -10262 7615 -10228 7649
rect -10262 7547 -10228 7581
rect -10262 7479 -10228 7513
rect -10478 7412 -10444 7446
rect -10086 7955 -10052 7989
rect -10086 7887 -10052 7921
rect -10086 7819 -10052 7853
rect -10086 7751 -10052 7785
rect -10086 7683 -10052 7717
rect -10086 7615 -10052 7649
rect -10086 7547 -10052 7581
rect -10086 7479 -10052 7513
rect -9910 7955 -9876 7989
rect -9662 7953 -9628 7987
rect -9910 7887 -9876 7921
rect -9910 7819 -9876 7853
rect -9910 7751 -9876 7785
rect -9910 7683 -9876 7717
rect -9910 7615 -9876 7649
rect -9910 7547 -9876 7581
rect -9910 7479 -9876 7513
rect -9662 7497 -9628 7531
rect -9662 7041 -9628 7075
rect -10604 6572 -10570 6606
rect -10604 6504 -10570 6538
rect -10604 6436 -10570 6470
rect -9748 6572 -9714 6606
rect -9748 6504 -9714 6538
rect -9748 6436 -9714 6470
rect -8092 6572 -8058 6606
rect -8092 6504 -8058 6538
rect -8092 6436 -8058 6470
rect -6436 6572 -6402 6606
rect -6436 6504 -6402 6538
rect -6436 6436 -6402 6470
rect -5580 6572 -5546 6606
rect -5580 6504 -5546 6538
rect -5580 6436 -5546 6470
rect -10339 6112 -10305 6146
rect -10339 6044 -10305 6078
rect -10339 5976 -10305 6010
rect -10163 6112 -10129 6146
rect -10163 6044 -10129 6078
rect -10163 5976 -10129 6010
<< mvpdiffc >>
rect 5776 12513 5810 12547
rect 5776 12445 5810 12479
rect 5952 12513 5986 12547
rect 5952 12445 5986 12479
rect 6134 12513 6168 12547
rect 6134 12445 6168 12479
rect 6310 12513 6344 12547
rect 6310 12445 6344 12479
rect 5860 12190 5894 12224
rect 5928 12190 5962 12224
rect 5996 12190 6030 12224
rect 6064 12190 6098 12224
rect 6132 12190 6166 12224
rect 6200 12190 6234 12224
rect 6268 12190 6302 12224
rect 6336 12190 6370 12224
rect 5860 12014 5894 12048
rect 5928 12014 5962 12048
rect 5996 12014 6030 12048
rect 6064 12014 6098 12048
rect 6132 12014 6166 12048
rect 6200 12014 6234 12048
rect 6268 12014 6302 12048
rect 6336 12014 6370 12048
rect 5860 11838 5894 11872
rect 5928 11838 5962 11872
rect 5996 11838 6030 11872
rect 6064 11838 6098 11872
rect 6132 11838 6166 11872
rect 6200 11838 6234 11872
rect 6268 11838 6302 11872
rect 6336 11838 6370 11872
rect 5860 11662 5894 11696
rect 5928 11662 5962 11696
rect 5996 11662 6030 11696
rect 6064 11662 6098 11696
rect 6132 11662 6166 11696
rect 6200 11662 6234 11696
rect 6268 11662 6302 11696
rect 6336 11662 6370 11696
rect 5860 11406 5894 11440
rect 5928 11406 5962 11440
rect 5996 11406 6030 11440
rect 6064 11406 6098 11440
rect 6132 11406 6166 11440
rect 6200 11406 6234 11440
rect 6268 11406 6302 11440
rect 6336 11406 6370 11440
rect 5860 11150 5894 11184
rect 5928 11150 5962 11184
rect 5996 11150 6030 11184
rect 6064 11150 6098 11184
rect 6132 11150 6166 11184
rect 6200 11150 6234 11184
rect 6268 11150 6302 11184
rect 6336 11150 6370 11184
rect 5860 10894 5894 10928
rect 5928 10894 5962 10928
rect 5996 10894 6030 10928
rect 6064 10894 6098 10928
rect 6132 10894 6166 10928
rect 6200 10894 6234 10928
rect 6268 10894 6302 10928
rect 6336 10894 6370 10928
rect 5860 10638 5894 10672
rect 5928 10638 5962 10672
rect 5996 10638 6030 10672
rect 6064 10638 6098 10672
rect 6132 10638 6166 10672
rect 6200 10638 6234 10672
rect 6268 10638 6302 10672
rect 6336 10638 6370 10672
rect 5860 10382 5894 10416
rect 5928 10382 5962 10416
rect 5996 10382 6030 10416
rect 6064 10382 6098 10416
rect 6132 10382 6166 10416
rect 6200 10382 6234 10416
rect 6268 10382 6302 10416
rect 6336 10382 6370 10416
rect 5860 10126 5894 10160
rect 5928 10126 5962 10160
rect 5996 10126 6030 10160
rect 6064 10126 6098 10160
rect 6132 10126 6166 10160
rect 6200 10126 6234 10160
rect 6268 10126 6302 10160
rect 6336 10126 6370 10160
rect 5860 9870 5894 9904
rect 5928 9870 5962 9904
rect 5996 9870 6030 9904
rect 6064 9870 6098 9904
rect 6132 9870 6166 9904
rect 6200 9870 6234 9904
rect 6268 9870 6302 9904
rect 6336 9870 6370 9904
rect 5860 9614 5894 9648
rect 5928 9614 5962 9648
rect 5996 9614 6030 9648
rect 6064 9614 6098 9648
rect 6132 9614 6166 9648
rect 6200 9614 6234 9648
rect 6268 9614 6302 9648
rect 6336 9614 6370 9648
rect 5913 9386 5947 9420
rect 5913 9318 5947 9352
rect 5913 9250 5947 9284
rect 6089 9386 6123 9420
rect 6089 9318 6123 9352
rect 6089 9250 6123 9284
rect 6265 9386 6299 9420
rect 6265 9318 6299 9352
rect 6265 9250 6299 9284
<< psubdiff >>
rect -10466 7122 -10432 7156
rect -10398 7122 -10358 7156
rect -10324 7122 -10284 7156
rect -10250 7122 -10210 7156
rect -10176 7122 -10135 7156
rect -10101 7122 -10060 7156
rect -10026 7122 -9985 7156
rect -9951 7122 -9910 7156
rect -9876 7122 -9842 7156
rect -10466 7088 -9842 7122
rect -10466 7054 -10432 7088
rect -10398 7054 -10358 7088
rect -10324 7054 -10284 7088
rect -10250 7054 -10210 7088
rect -10176 7054 -10135 7088
rect -10101 7054 -10060 7088
rect -10026 7054 -9985 7088
rect -9951 7054 -9910 7088
rect -9876 7054 -9842 7088
rect -10466 7020 -9842 7054
rect -10466 6986 -10432 7020
rect -10398 6986 -10358 7020
rect -10324 6986 -10284 7020
rect -10250 6986 -10210 7020
rect -10176 6986 -10135 7020
rect -10101 6986 -10060 7020
rect -10026 6986 -9985 7020
rect -9951 6986 -9910 7020
rect -9876 6986 -9842 7020
rect -10466 6952 -9842 6986
rect -10466 6918 -10432 6952
rect -10398 6918 -10358 6952
rect -10324 6918 -10284 6952
rect -10250 6918 -10210 6952
rect -10176 6918 -10135 6952
rect -10101 6918 -10060 6952
rect -10026 6918 -9985 6952
rect -9951 6918 -9910 6952
rect -9876 6918 -9842 6952
rect -10466 6884 -9842 6918
rect -10466 6850 -10432 6884
rect -10398 6850 -10358 6884
rect -10324 6850 -10284 6884
rect -10250 6850 -10210 6884
rect -10176 6850 -10135 6884
rect -10101 6850 -10060 6884
rect -10026 6850 -9985 6884
rect -9951 6850 -9910 6884
rect -9876 6850 -9842 6884
rect -10466 6798 -9842 6850
rect -10466 6696 -10442 6798
rect -2792 6764 -2757 6798
rect -2723 6764 -2688 6798
rect -2654 6764 -2619 6798
rect -2585 6764 -2550 6798
rect -2516 6764 -2481 6798
rect -2447 6764 -2412 6798
rect -2378 6764 -2343 6798
rect -2309 6764 -2274 6798
rect -2240 6764 -2205 6798
rect -2171 6764 -2136 6798
rect -2102 6764 -2067 6798
rect -2033 6764 -1998 6798
rect -1964 6764 -1929 6798
rect -1895 6764 -1871 6798
rect -2792 6730 -1871 6764
rect -2792 6696 -2757 6730
rect -2723 6696 -2688 6730
rect -2654 6696 -2619 6730
rect -2585 6696 -2550 6730
rect -2516 6696 -2481 6730
rect -2447 6696 -2412 6730
rect -2378 6696 -2343 6730
rect -2309 6696 -2274 6730
rect -2240 6696 -2205 6730
rect -2171 6696 -2136 6730
rect -2102 6696 -2067 6730
rect -2033 6696 -1998 6730
rect -1964 6696 -1929 6730
rect -1895 6696 -1871 6730
<< psubdiffcont >>
rect -10432 7122 -10398 7156
rect -10358 7122 -10324 7156
rect -10284 7122 -10250 7156
rect -10210 7122 -10176 7156
rect -10135 7122 -10101 7156
rect -10060 7122 -10026 7156
rect -9985 7122 -9951 7156
rect -9910 7122 -9876 7156
rect -10432 7054 -10398 7088
rect -10358 7054 -10324 7088
rect -10284 7054 -10250 7088
rect -10210 7054 -10176 7088
rect -10135 7054 -10101 7088
rect -10060 7054 -10026 7088
rect -9985 7054 -9951 7088
rect -9910 7054 -9876 7088
rect -10432 6986 -10398 7020
rect -10358 6986 -10324 7020
rect -10284 6986 -10250 7020
rect -10210 6986 -10176 7020
rect -10135 6986 -10101 7020
rect -10060 6986 -10026 7020
rect -9985 6986 -9951 7020
rect -9910 6986 -9876 7020
rect -10432 6918 -10398 6952
rect -10358 6918 -10324 6952
rect -10284 6918 -10250 6952
rect -10210 6918 -10176 6952
rect -10135 6918 -10101 6952
rect -10060 6918 -10026 6952
rect -9985 6918 -9951 6952
rect -9910 6918 -9876 6952
rect -10432 6850 -10398 6884
rect -10358 6850 -10324 6884
rect -10284 6850 -10250 6884
rect -10210 6850 -10176 6884
rect -10135 6850 -10101 6884
rect -10060 6850 -10026 6884
rect -9985 6850 -9951 6884
rect -9910 6850 -9876 6884
rect -10442 6696 -2792 6798
rect -2757 6764 -2723 6798
rect -2688 6764 -2654 6798
rect -2619 6764 -2585 6798
rect -2550 6764 -2516 6798
rect -2481 6764 -2447 6798
rect -2412 6764 -2378 6798
rect -2343 6764 -2309 6798
rect -2274 6764 -2240 6798
rect -2205 6764 -2171 6798
rect -2136 6764 -2102 6798
rect -2067 6764 -2033 6798
rect -1998 6764 -1964 6798
rect -1929 6764 -1895 6798
rect -2757 6696 -2723 6730
rect -2688 6696 -2654 6730
rect -2619 6696 -2585 6730
rect -2550 6696 -2516 6730
rect -2481 6696 -2447 6730
rect -2412 6696 -2378 6730
rect -2343 6696 -2309 6730
rect -2274 6696 -2240 6730
rect -2205 6696 -2171 6730
rect -2136 6696 -2102 6730
rect -2067 6696 -2033 6730
rect -1998 6696 -1964 6730
rect -1929 6696 -1895 6730
<< poly >>
rect 5807 12655 5941 12671
rect 5807 12621 5823 12655
rect 5857 12621 5891 12655
rect 5925 12621 5941 12655
rect 5807 12605 5941 12621
rect 6165 12655 6299 12671
rect 6165 12621 6181 12655
rect 6215 12621 6249 12655
rect 6283 12621 6299 12655
rect 6165 12605 6299 12621
rect 5821 12573 5941 12605
rect 6179 12573 6299 12605
rect 5821 12401 5941 12433
rect 6179 12401 6299 12433
rect 5684 12179 5750 12193
rect 5684 12177 5782 12179
rect 5684 12143 5700 12177
rect 5734 12143 5782 12177
rect 5684 12109 5782 12143
rect 5684 12075 5700 12109
rect 5734 12075 5782 12109
rect 5684 12059 5782 12075
rect 6382 12059 6414 12179
rect 5684 11987 5782 12003
rect 5684 11953 5700 11987
rect 5734 11953 5782 11987
rect 5684 11911 5782 11953
rect 5684 11877 5700 11911
rect 5734 11883 5782 11911
rect 6382 11883 6414 12003
rect 5734 11877 5750 11883
rect 5684 11834 5750 11877
rect 5684 11800 5700 11834
rect 5734 11827 5750 11834
rect 5734 11800 5782 11827
rect 5684 11757 5782 11800
rect 5684 11723 5700 11757
rect 5734 11723 5782 11757
rect 5684 11707 5782 11723
rect 6382 11707 6414 11827
rect 5684 11635 5782 11651
rect 5684 11601 5700 11635
rect 5734 11601 5782 11635
rect 5684 11557 5782 11601
rect 5684 11523 5700 11557
rect 5734 11523 5782 11557
rect 5684 11479 5782 11523
rect 5684 11445 5700 11479
rect 5734 11451 5782 11479
rect 6382 11451 6414 11651
rect 5734 11445 5750 11451
rect 5684 11401 5750 11445
rect 5684 11367 5700 11401
rect 5734 11395 5750 11401
rect 5734 11367 5782 11395
rect 5684 11323 5782 11367
rect 5684 11289 5700 11323
rect 5734 11289 5782 11323
rect 5684 11245 5782 11289
rect 5684 11211 5700 11245
rect 5734 11211 5782 11245
rect 5684 11195 5782 11211
rect 6382 11195 6414 11395
rect 5684 11123 5782 11139
rect 5684 11089 5700 11123
rect 5734 11089 5782 11123
rect 5684 11045 5782 11089
rect 5684 11011 5700 11045
rect 5734 11011 5782 11045
rect 5684 10967 5782 11011
rect 5684 10933 5700 10967
rect 5734 10939 5782 10967
rect 6382 10939 6414 11139
rect 5734 10933 5750 10939
rect 5684 10889 5750 10933
rect 5684 10855 5700 10889
rect 5734 10883 5750 10889
rect 5734 10855 5782 10883
rect 5684 10811 5782 10855
rect 5684 10777 5700 10811
rect 5734 10777 5782 10811
rect 5684 10733 5782 10777
rect 5684 10699 5700 10733
rect 5734 10699 5782 10733
rect 5684 10683 5782 10699
rect 6382 10683 6414 10883
rect 5684 10611 5782 10627
rect 5684 10577 5700 10611
rect 5734 10577 5782 10611
rect 5684 10533 5782 10577
rect 5684 10499 5700 10533
rect 5734 10499 5782 10533
rect 5684 10455 5782 10499
rect 5684 10421 5700 10455
rect 5734 10427 5782 10455
rect 6382 10427 6414 10627
rect 5734 10421 5750 10427
rect 5684 10377 5750 10421
rect 5684 10343 5700 10377
rect 5734 10371 5750 10377
rect 5734 10343 5782 10371
rect 5684 10299 5782 10343
rect 5684 10265 5700 10299
rect 5734 10265 5782 10299
rect 5684 10221 5782 10265
rect 5684 10187 5700 10221
rect 5734 10187 5782 10221
rect 5684 10171 5782 10187
rect 6382 10171 6414 10371
rect 5684 10099 5782 10115
rect 5684 10065 5700 10099
rect 5734 10065 5782 10099
rect 5684 10021 5782 10065
rect 5684 9987 5700 10021
rect 5734 9987 5782 10021
rect 5684 9943 5782 9987
rect 5684 9909 5700 9943
rect 5734 9915 5782 9943
rect 6382 9915 6414 10115
rect 5734 9909 5750 9915
rect 5684 9865 5750 9909
rect 5684 9831 5700 9865
rect 5734 9859 5750 9865
rect 5734 9831 5782 9859
rect 5684 9787 5782 9831
rect 5684 9753 5700 9787
rect 5734 9753 5782 9787
rect 5684 9709 5782 9753
rect 5684 9675 5700 9709
rect 5734 9675 5782 9709
rect 5684 9659 5782 9675
rect 6382 9659 6414 9859
rect 5958 9432 6078 9464
rect 6134 9432 6254 9464
rect 5958 9200 6078 9232
rect 6134 9200 6254 9232
rect 5958 9184 6254 9200
rect 5958 9150 5974 9184
rect 6008 9150 6050 9184
rect 6084 9150 6127 9184
rect 6161 9150 6204 9184
rect 6238 9150 6254 9184
rect 5958 9134 6254 9150
rect -10217 8001 -10097 8033
rect -10041 8001 -9921 8033
rect -10548 7457 -10516 7857
rect -10432 7841 -10334 7857
rect -10432 7807 -10384 7841
rect -10350 7807 -10334 7841
rect -10432 7757 -10334 7807
rect -10432 7723 -10384 7757
rect -10350 7723 -10334 7757
rect -10432 7673 -10334 7723
rect -10432 7639 -10384 7673
rect -10350 7639 -10334 7673
rect -10432 7590 -10334 7639
rect -10432 7556 -10384 7590
rect -10350 7556 -10334 7590
rect -10432 7507 -10334 7556
rect -10432 7473 -10384 7507
rect -10350 7473 -10334 7507
rect -10432 7457 -10334 7473
rect -9732 7542 -9700 7942
rect -9616 7926 -9518 7942
rect -9616 7892 -9568 7926
rect -9534 7892 -9518 7926
rect -9616 7854 -9518 7892
rect -9616 7820 -9568 7854
rect -9534 7820 -9518 7854
rect -9616 7782 -9518 7820
rect -9616 7748 -9568 7782
rect -9534 7748 -9518 7782
rect -9616 7710 -9518 7748
rect -9616 7676 -9568 7710
rect -9534 7676 -9518 7710
rect -9616 7638 -9518 7676
rect -9616 7604 -9568 7638
rect -9534 7604 -9518 7638
rect -9616 7566 -9518 7604
rect -9616 7542 -9568 7566
rect -9584 7532 -9568 7542
rect -9534 7532 -9518 7566
rect -9584 7494 -9518 7532
rect -9584 7486 -9568 7494
rect -10217 7369 -10097 7401
rect -10231 7353 -10097 7369
rect -10231 7319 -10215 7353
rect -10181 7319 -10147 7353
rect -10113 7319 -10097 7353
rect -10231 7303 -10097 7319
rect -10041 7369 -9921 7401
rect -10041 7353 -9907 7369
rect -10041 7319 -10025 7353
rect -9991 7319 -9957 7353
rect -9923 7319 -9907 7353
rect -10041 7303 -9907 7319
rect -9732 7086 -9700 7486
rect -9616 7460 -9568 7486
rect -9534 7460 -9518 7494
rect -9616 7422 -9518 7460
rect -9616 7388 -9568 7422
rect -9534 7388 -9518 7422
rect -9616 7350 -9518 7388
rect -9616 7316 -9568 7350
rect -9534 7316 -9518 7350
rect -9616 7278 -9518 7316
rect -9616 7244 -9568 7278
rect -9534 7244 -9518 7278
rect -9616 7207 -9518 7244
rect -9616 7173 -9568 7207
rect -9534 7173 -9518 7207
rect -9616 7136 -9518 7173
rect -9616 7102 -9568 7136
rect -9534 7102 -9518 7136
rect -9616 7086 -9518 7102
rect -10559 6618 -9759 6650
rect -9703 6618 -8103 6650
rect -8047 6618 -6447 6650
rect -6391 6618 -5591 6650
rect -10559 6370 -9759 6418
rect -10559 6336 -10543 6370
rect -10509 6336 -10470 6370
rect -10436 6336 -10397 6370
rect -10363 6336 -10324 6370
rect -10290 6336 -10251 6370
rect -10217 6336 -10178 6370
rect -10144 6336 -10105 6370
rect -10071 6336 -10031 6370
rect -9997 6336 -9957 6370
rect -9923 6336 -9883 6370
rect -9849 6336 -9809 6370
rect -9775 6336 -9759 6370
rect -10559 6320 -9759 6336
rect -9703 6370 -8103 6418
rect -9703 6336 -9687 6370
rect -9653 6336 -9618 6370
rect -9584 6336 -9549 6370
rect -9515 6336 -9480 6370
rect -9446 6336 -9411 6370
rect -9377 6336 -9342 6370
rect -9308 6336 -9273 6370
rect -9239 6336 -9203 6370
rect -9169 6336 -9133 6370
rect -9099 6336 -9063 6370
rect -9029 6336 -8993 6370
rect -8959 6336 -8923 6370
rect -8889 6336 -8853 6370
rect -8819 6336 -8783 6370
rect -8749 6336 -8713 6370
rect -8679 6336 -8643 6370
rect -8609 6336 -8573 6370
rect -8539 6336 -8503 6370
rect -8469 6336 -8433 6370
rect -8399 6336 -8363 6370
rect -8329 6336 -8293 6370
rect -8259 6336 -8223 6370
rect -8189 6336 -8153 6370
rect -8119 6336 -8103 6370
rect -9703 6320 -8103 6336
rect -8047 6370 -6447 6418
rect -8047 6336 -8031 6370
rect -7997 6336 -7962 6370
rect -7928 6336 -7893 6370
rect -7859 6336 -7824 6370
rect -7790 6336 -7755 6370
rect -7721 6336 -7686 6370
rect -7652 6336 -7617 6370
rect -7583 6336 -7547 6370
rect -7513 6336 -7477 6370
rect -7443 6336 -7407 6370
rect -7373 6336 -7337 6370
rect -7303 6336 -7267 6370
rect -7233 6336 -7197 6370
rect -7163 6336 -7127 6370
rect -7093 6336 -7057 6370
rect -7023 6336 -6987 6370
rect -6953 6336 -6917 6370
rect -6883 6336 -6847 6370
rect -6813 6336 -6777 6370
rect -6743 6336 -6707 6370
rect -6673 6336 -6637 6370
rect -6603 6336 -6567 6370
rect -6533 6336 -6497 6370
rect -6463 6336 -6447 6370
rect -8047 6320 -6447 6336
rect -6391 6370 -5591 6418
rect -6391 6336 -6375 6370
rect -6341 6336 -6302 6370
rect -6268 6336 -6229 6370
rect -6195 6336 -6156 6370
rect -6122 6336 -6083 6370
rect -6049 6336 -6010 6370
rect -5976 6336 -5937 6370
rect -5903 6336 -5863 6370
rect -5829 6336 -5789 6370
rect -5755 6336 -5715 6370
rect -5681 6336 -5641 6370
rect -5607 6336 -5591 6370
rect -6391 6320 -5591 6336
rect -10294 6246 -10160 6262
rect -10294 6212 -10278 6246
rect -10244 6212 -10210 6246
rect -10176 6212 -10160 6246
rect -10294 6196 -10160 6212
rect -10294 6164 -10174 6196
rect -10294 5932 -10174 5964
<< polycont >>
rect 5823 12621 5857 12655
rect 5891 12621 5925 12655
rect 6181 12621 6215 12655
rect 6249 12621 6283 12655
rect 5700 12143 5734 12177
rect 5700 12075 5734 12109
rect 5700 11953 5734 11987
rect 5700 11877 5734 11911
rect 5700 11800 5734 11834
rect 5700 11723 5734 11757
rect 5700 11601 5734 11635
rect 5700 11523 5734 11557
rect 5700 11445 5734 11479
rect 5700 11367 5734 11401
rect 5700 11289 5734 11323
rect 5700 11211 5734 11245
rect 5700 11089 5734 11123
rect 5700 11011 5734 11045
rect 5700 10933 5734 10967
rect 5700 10855 5734 10889
rect 5700 10777 5734 10811
rect 5700 10699 5734 10733
rect 5700 10577 5734 10611
rect 5700 10499 5734 10533
rect 5700 10421 5734 10455
rect 5700 10343 5734 10377
rect 5700 10265 5734 10299
rect 5700 10187 5734 10221
rect 5700 10065 5734 10099
rect 5700 9987 5734 10021
rect 5700 9909 5734 9943
rect 5700 9831 5734 9865
rect 5700 9753 5734 9787
rect 5700 9675 5734 9709
rect 5974 9150 6008 9184
rect 6050 9150 6084 9184
rect 6127 9150 6161 9184
rect 6204 9150 6238 9184
rect -10384 7807 -10350 7841
rect -10384 7723 -10350 7757
rect -10384 7639 -10350 7673
rect -10384 7556 -10350 7590
rect -10384 7473 -10350 7507
rect -9568 7892 -9534 7926
rect -9568 7820 -9534 7854
rect -9568 7748 -9534 7782
rect -9568 7676 -9534 7710
rect -9568 7604 -9534 7638
rect -9568 7532 -9534 7566
rect -10215 7319 -10181 7353
rect -10147 7319 -10113 7353
rect -10025 7319 -9991 7353
rect -9957 7319 -9923 7353
rect -9568 7460 -9534 7494
rect -9568 7388 -9534 7422
rect -9568 7316 -9534 7350
rect -9568 7244 -9534 7278
rect -9568 7173 -9534 7207
rect -9568 7102 -9534 7136
rect -10543 6336 -10509 6370
rect -10470 6336 -10436 6370
rect -10397 6336 -10363 6370
rect -10324 6336 -10290 6370
rect -10251 6336 -10217 6370
rect -10178 6336 -10144 6370
rect -10105 6336 -10071 6370
rect -10031 6336 -9997 6370
rect -9957 6336 -9923 6370
rect -9883 6336 -9849 6370
rect -9809 6336 -9775 6370
rect -9687 6336 -9653 6370
rect -9618 6336 -9584 6370
rect -9549 6336 -9515 6370
rect -9480 6336 -9446 6370
rect -9411 6336 -9377 6370
rect -9342 6336 -9308 6370
rect -9273 6336 -9239 6370
rect -9203 6336 -9169 6370
rect -9133 6336 -9099 6370
rect -9063 6336 -9029 6370
rect -8993 6336 -8959 6370
rect -8923 6336 -8889 6370
rect -8853 6336 -8819 6370
rect -8783 6336 -8749 6370
rect -8713 6336 -8679 6370
rect -8643 6336 -8609 6370
rect -8573 6336 -8539 6370
rect -8503 6336 -8469 6370
rect -8433 6336 -8399 6370
rect -8363 6336 -8329 6370
rect -8293 6336 -8259 6370
rect -8223 6336 -8189 6370
rect -8153 6336 -8119 6370
rect -8031 6336 -7997 6370
rect -7962 6336 -7928 6370
rect -7893 6336 -7859 6370
rect -7824 6336 -7790 6370
rect -7755 6336 -7721 6370
rect -7686 6336 -7652 6370
rect -7617 6336 -7583 6370
rect -7547 6336 -7513 6370
rect -7477 6336 -7443 6370
rect -7407 6336 -7373 6370
rect -7337 6336 -7303 6370
rect -7267 6336 -7233 6370
rect -7197 6336 -7163 6370
rect -7127 6336 -7093 6370
rect -7057 6336 -7023 6370
rect -6987 6336 -6953 6370
rect -6917 6336 -6883 6370
rect -6847 6336 -6813 6370
rect -6777 6336 -6743 6370
rect -6707 6336 -6673 6370
rect -6637 6336 -6603 6370
rect -6567 6336 -6533 6370
rect -6497 6336 -6463 6370
rect -6375 6336 -6341 6370
rect -6302 6336 -6268 6370
rect -6229 6336 -6195 6370
rect -6156 6336 -6122 6370
rect -6083 6336 -6049 6370
rect -6010 6336 -5976 6370
rect -5937 6336 -5903 6370
rect -5863 6336 -5829 6370
rect -5789 6336 -5755 6370
rect -5715 6336 -5681 6370
rect -5641 6336 -5607 6370
rect -10278 6212 -10244 6246
rect -10210 6212 -10176 6246
<< locali >>
rect 6112 12672 6299 12706
rect 6078 12655 6299 12672
rect 5807 12621 5823 12655
rect 5857 12621 5891 12655
rect 5929 12621 5941 12655
rect 6078 12634 6181 12655
rect 6112 12621 6181 12634
rect 6215 12621 6249 12655
rect 6283 12621 6299 12655
rect 5953 12563 6168 12564
rect 5776 12547 5810 12563
rect 5776 12479 5810 12509
rect 5776 12429 5810 12437
rect 5952 12547 6168 12563
rect 5986 12543 6134 12547
rect 5992 12513 6134 12543
rect 5952 12509 5958 12513
rect 5992 12509 6168 12513
rect 5952 12479 6168 12509
rect 5986 12471 6134 12479
rect 5992 12445 6134 12471
rect 5952 12437 5958 12445
rect 5992 12437 6168 12445
rect 5952 12429 6168 12437
rect 6310 12547 6344 12563
rect 6310 12479 6348 12513
rect 6344 12475 6348 12479
rect 6310 12441 6314 12445
rect 6310 12429 6344 12441
rect 5953 12425 6168 12429
rect 5562 12303 6387 12337
rect 5528 12265 6387 12303
rect 5562 12236 6387 12265
rect 5844 12224 6387 12236
rect 5700 12177 5734 12193
rect 5844 12190 5860 12224
rect 5894 12190 5928 12224
rect 5962 12190 5996 12224
rect 6030 12190 6064 12224
rect 6098 12190 6132 12224
rect 6166 12190 6200 12224
rect 6234 12190 6268 12224
rect 6302 12190 6336 12224
rect 6370 12193 6387 12224
rect 6370 12190 6386 12193
rect 5700 12109 5734 12143
rect 5700 12059 5734 12071
rect 5844 12014 5856 12048
rect 5894 12014 5928 12048
rect 5962 12014 5986 12048
rect 6030 12014 6064 12048
rect 6098 12014 6132 12048
rect 6166 12014 6200 12048
rect 6234 12014 6268 12048
rect 6302 12014 6336 12048
rect 6370 12014 6386 12048
rect 5700 11991 5734 12003
rect 5700 11912 5734 11953
rect 5700 11834 5734 11877
rect 5844 11838 5860 11872
rect 5894 11838 5928 11872
rect 5962 11838 5996 11872
rect 6030 11838 6064 11872
rect 6098 11838 6132 11872
rect 6166 11838 6200 11872
rect 6234 11838 6268 11872
rect 6302 11838 6336 11872
rect 6370 11838 6386 11872
rect 6248 11834 6282 11838
rect 5700 11757 5734 11799
rect 5700 11707 5734 11719
rect 5844 11662 5856 11696
rect 5894 11662 5928 11696
rect 5962 11662 5986 11696
rect 6030 11662 6064 11696
rect 6098 11662 6132 11696
rect 6166 11662 6200 11696
rect 6234 11662 6268 11696
rect 6302 11662 6336 11696
rect 6370 11662 6386 11696
rect 5700 11639 5734 11651
rect 5700 11560 5734 11601
rect 5700 11481 5734 11523
rect 5700 11401 5734 11445
rect 5845 11442 6163 11476
rect 6197 11442 6386 11476
rect 5845 11440 6386 11442
rect 5844 11406 5860 11440
rect 5894 11406 5928 11440
rect 5962 11406 5996 11440
rect 6030 11406 6064 11440
rect 6098 11406 6132 11440
rect 6166 11406 6200 11440
rect 6234 11406 6268 11440
rect 6302 11406 6336 11440
rect 6370 11406 6386 11440
rect 5845 11401 6386 11406
rect 5845 11367 6163 11401
rect 6197 11367 6386 11401
rect 5700 11323 5734 11367
rect 5700 11245 5734 11287
rect 5700 11195 5734 11207
rect 5844 11150 5856 11184
rect 5894 11150 5928 11184
rect 5962 11150 5986 11184
rect 6030 11150 6064 11184
rect 6098 11150 6132 11184
rect 6166 11150 6200 11184
rect 6234 11150 6268 11184
rect 6302 11150 6336 11184
rect 6370 11150 6386 11184
rect 5700 11127 5734 11139
rect 5700 11048 5734 11089
rect 5700 10969 5734 11011
rect 5700 10889 5734 10933
rect 5845 10930 6163 10964
rect 6197 10930 6386 10964
rect 5845 10928 6386 10930
rect 5844 10894 5860 10928
rect 5894 10894 5928 10928
rect 5962 10894 5996 10928
rect 6030 10894 6064 10928
rect 6098 10894 6132 10928
rect 6166 10894 6200 10928
rect 6234 10894 6268 10928
rect 6302 10894 6336 10928
rect 6370 10894 6386 10928
rect 5845 10889 6386 10894
rect 5845 10855 6163 10889
rect 6197 10855 6386 10889
rect 5700 10811 5734 10855
rect 5700 10733 5734 10775
rect 5700 10683 5734 10695
rect 5844 10638 5856 10672
rect 5894 10638 5928 10672
rect 5962 10638 5986 10672
rect 6030 10638 6064 10672
rect 6098 10638 6132 10672
rect 6166 10638 6200 10672
rect 6234 10638 6268 10672
rect 6302 10638 6336 10672
rect 6370 10638 6386 10672
rect 5700 10615 5734 10627
rect 5700 10536 5734 10577
rect 5700 10457 5734 10499
rect 5700 10377 5734 10421
rect 5845 10417 6078 10451
rect 6112 10417 6386 10451
rect 5845 10416 6386 10417
rect 5844 10382 5860 10416
rect 5894 10382 5928 10416
rect 5962 10382 5996 10416
rect 6030 10382 6064 10416
rect 6098 10382 6132 10416
rect 6166 10382 6200 10416
rect 6234 10382 6268 10416
rect 6302 10382 6336 10416
rect 6370 10382 6386 10416
rect 5700 10299 5734 10343
rect 5845 10376 6386 10382
rect 5845 10342 6078 10376
rect 6112 10342 6386 10376
rect 5700 10221 5734 10263
rect 5700 10171 5734 10183
rect 5844 10126 5856 10160
rect 5894 10126 5928 10160
rect 5962 10126 5986 10160
rect 6030 10126 6064 10160
rect 6098 10126 6132 10160
rect 6166 10126 6200 10160
rect 6234 10126 6268 10160
rect 6302 10126 6336 10160
rect 6370 10126 6386 10160
rect 5700 10103 5734 10115
rect 5700 10024 5734 10065
rect 5700 9945 5734 9987
rect 5700 9865 5734 9909
rect 5845 9905 6078 9939
rect 6112 9905 6386 9939
rect 5845 9904 6386 9905
rect 5844 9870 5860 9904
rect 5894 9870 5928 9904
rect 5962 9870 5996 9904
rect 6030 9870 6064 9904
rect 6098 9870 6132 9904
rect 6166 9870 6200 9904
rect 6234 9870 6268 9904
rect 6302 9870 6336 9904
rect 6370 9870 6386 9904
rect 5700 9787 5734 9831
rect 5845 9864 6386 9870
rect 5845 9830 6078 9864
rect 6112 9830 6386 9864
rect 5700 9709 5734 9751
rect 5700 9659 5734 9671
rect 5844 9614 5856 9648
rect 5894 9614 5928 9648
rect 5962 9614 5986 9648
rect 6030 9614 6064 9648
rect 6098 9614 6132 9648
rect 6166 9614 6200 9648
rect 6234 9614 6268 9648
rect 6302 9614 6336 9648
rect 6370 9614 6386 9648
rect 5732 9566 5772 9568
rect 5806 9566 5812 9568
rect 5732 9528 5812 9566
rect 5732 9494 5772 9528
rect 5806 9494 5812 9528
rect 5732 9184 5812 9494
rect 5847 9471 6320 9560
rect 5847 9420 5947 9471
rect 6089 9423 6123 9436
rect 5847 9374 5913 9420
rect 5847 9352 5947 9374
rect 5847 9318 5913 9352
rect 5847 9284 5947 9318
rect 5847 9244 5913 9284
rect 6109 9420 6123 9423
rect 6075 9386 6089 9389
rect 6075 9352 6123 9386
rect 6075 9318 6089 9352
rect 6075 9302 6123 9318
rect 6109 9284 6123 9302
rect 5847 9234 5947 9244
rect 6089 9234 6123 9250
rect 6264 9420 6320 9471
rect 6264 9386 6265 9420
rect 6299 9386 6320 9420
rect 6264 9352 6320 9386
rect 6264 9318 6265 9352
rect 6299 9318 6320 9352
rect 6264 9284 6320 9318
rect 6264 9250 6265 9284
rect 6299 9250 6320 9284
rect 6264 9234 6320 9250
rect 5732 9178 5974 9184
rect 6008 9178 6050 9184
rect 5732 9144 5969 9178
rect 6008 9150 6043 9178
rect 6084 9150 6127 9184
rect 6161 9150 6204 9184
rect 6238 9150 6282 9184
rect 6003 9144 6043 9150
rect 6077 9144 6282 9150
rect 5732 9085 6282 9144
rect 5606 9049 5640 9072
rect 6333 9049 6367 9072
rect 5606 9034 6367 9049
rect 5640 9000 6333 9034
rect 5606 8988 6367 9000
rect 5706 8906 5778 8940
rect 5812 8917 6283 8940
rect 5812 8906 6249 8917
rect 5706 8883 6249 8906
rect 5706 8879 6283 8883
rect 5778 8868 5812 8879
rect 6249 8844 6283 8879
rect -10262 7989 -10228 8005
rect -10262 7921 -10228 7955
rect -10500 7902 -10462 7908
rect -10500 7874 -10478 7902
rect -10494 7868 -10478 7874
rect -10444 7868 -10428 7874
rect -10382 7857 -10348 7859
rect -10384 7841 -10348 7857
rect -10350 7808 -10348 7841
rect -10384 7774 -10382 7807
rect -10384 7757 -10348 7774
rect -10350 7723 -10348 7757
rect -10384 7689 -10382 7723
rect -10384 7673 -10348 7689
rect -10350 7639 -10348 7673
rect -10384 7638 -10348 7639
rect -10384 7604 -10382 7638
rect -10384 7590 -10348 7604
rect -10350 7556 -10348 7590
rect -10384 7553 -10348 7556
rect -10384 7519 -10382 7553
rect -10262 7853 -10228 7859
rect -10262 7808 -10228 7819
rect -10262 7723 -10228 7751
rect -10262 7649 -10228 7683
rect -10262 7581 -10228 7604
rect -10384 7507 -10350 7519
rect -10384 7457 -10350 7473
rect -10262 7513 -10228 7519
rect -10262 7463 -10228 7479
rect -10086 7989 -10052 8005
rect -10086 7921 -10052 7955
rect -10086 7853 -10052 7887
rect -10086 7785 -10052 7819
rect -10086 7717 -10052 7751
rect -10086 7670 -10052 7683
rect -10086 7589 -10052 7615
rect -10086 7513 -10052 7547
rect -10086 7463 -10052 7475
rect -9910 7993 -9876 8005
rect -9910 7921 -9876 7955
rect -9687 7953 -9662 7962
rect -9628 7953 -9612 7987
rect -9687 7924 -9653 7953
rect -9568 7930 -9534 7942
rect -9910 7853 -9876 7877
rect -9910 7785 -9876 7795
rect -9910 7746 -9876 7751
rect -9910 7663 -9876 7683
rect -9910 7581 -9876 7615
rect -9568 7854 -9534 7892
rect -9568 7782 -9534 7815
rect -9568 7710 -9534 7734
rect -9568 7638 -9534 7653
rect -9910 7513 -9876 7546
rect -9687 7531 -9653 7538
rect -9568 7566 -9534 7572
rect -9687 7500 -9662 7531
rect -9628 7497 -9612 7531
rect -9568 7525 -9534 7532
rect -10519 7421 -10490 7446
rect -10519 7412 -10478 7421
rect -10444 7412 -10428 7446
rect -10519 7383 -10428 7412
rect -10519 7349 -10490 7383
rect -10456 7349 -10428 7383
rect -9568 7444 -9534 7460
rect -9995 7353 -9957 7365
rect -9568 7363 -9534 7388
rect -10519 7156 -10428 7349
rect -10231 7319 -10219 7353
rect -10181 7319 -10147 7353
rect -10113 7319 -10097 7353
rect -10041 7331 -10029 7353
rect -10041 7319 -10025 7331
rect -9991 7319 -9957 7353
rect -9923 7319 -9907 7353
rect -9568 7278 -9534 7316
rect -9568 7207 -9534 7244
rect -10519 7122 -10432 7156
rect -10398 7122 -10358 7156
rect -10324 7122 -10284 7156
rect -10250 7122 -10210 7156
rect -10176 7122 -10135 7156
rect -10101 7122 -10060 7156
rect -10026 7122 -9985 7156
rect -9951 7122 -9910 7156
rect -9876 7122 -9842 7156
rect -10519 7088 -9842 7122
rect -10519 7054 -10432 7088
rect -10398 7054 -10358 7088
rect -10324 7054 -10284 7088
rect -10250 7054 -10210 7088
rect -10176 7054 -10135 7088
rect -10101 7054 -10060 7088
rect -10026 7054 -9985 7088
rect -9951 7054 -9910 7088
rect -9876 7075 -9842 7088
rect -9568 7136 -9534 7173
rect -9568 7086 -9534 7102
rect -9876 7054 -9662 7075
rect -10519 7041 -9662 7054
rect -9628 7041 -9611 7075
rect -10519 7020 -9611 7041
rect -10519 6986 -10432 7020
rect -10398 6986 -10358 7020
rect -10324 6986 -10284 7020
rect -10250 6986 -10210 7020
rect -10176 6986 -10135 7020
rect -10101 6986 -10060 7020
rect -10026 6986 -9985 7020
rect -9951 6986 -9910 7020
rect -9876 6986 -9611 7020
rect -10519 6952 -9611 6986
rect -10519 6918 -10432 6952
rect -10398 6918 -10358 6952
rect -10324 6918 -10284 6952
rect -10250 6918 -10210 6952
rect -10176 6918 -10135 6952
rect -10101 6918 -10060 6952
rect -10026 6918 -9985 6952
rect -9951 6918 -9910 6952
rect -9876 6918 -9611 6952
rect -10519 6884 -9611 6918
rect -10519 6850 -10432 6884
rect -10398 6850 -10358 6884
rect -10324 6850 -10284 6884
rect -10250 6850 -10210 6884
rect -10176 6850 -10135 6884
rect -10101 6850 -10060 6884
rect -10026 6850 -9985 6884
rect -9951 6850 -9910 6884
rect -9876 6850 -9611 6884
rect -10519 6798 -9611 6850
rect -10466 6748 -10442 6798
rect -2792 6764 -2757 6798
rect -2723 6764 -2688 6798
rect -2654 6764 -2619 6798
rect -2585 6764 -2550 6798
rect -2516 6764 -2481 6798
rect -2447 6764 -2412 6798
rect -2378 6764 -2343 6798
rect -2309 6764 -2274 6798
rect -2240 6764 -2205 6798
rect -2171 6764 -2136 6798
rect -2102 6764 -2067 6798
rect -2033 6764 -1998 6798
rect -1964 6764 -1929 6798
rect -1895 6764 -1871 6798
rect -2792 6748 -1871 6764
rect -10466 6714 -10447 6748
rect -2792 6714 -2783 6748
rect -2749 6730 -2710 6748
rect -2676 6730 -2637 6748
rect -2603 6730 -2564 6748
rect -2530 6730 -2491 6748
rect -2457 6730 -2418 6748
rect -2384 6730 -2345 6748
rect -2311 6730 -2272 6748
rect -2238 6730 -2199 6748
rect -2165 6730 -2126 6748
rect -2092 6730 -2053 6748
rect -2019 6730 -1980 6748
rect -1946 6730 -1907 6748
rect -2723 6714 -2710 6730
rect -2654 6714 -2637 6730
rect -2585 6714 -2564 6730
rect -2516 6714 -2491 6730
rect -2447 6714 -2418 6730
rect -2378 6714 -2345 6730
rect -10466 6696 -10442 6714
rect -2792 6696 -2757 6714
rect -2723 6696 -2688 6714
rect -2654 6696 -2619 6714
rect -2585 6696 -2550 6714
rect -2516 6696 -2481 6714
rect -2447 6696 -2412 6714
rect -2378 6696 -2343 6714
rect -2309 6696 -2274 6730
rect -2238 6714 -2205 6730
rect -2165 6714 -2136 6730
rect -2092 6714 -2067 6730
rect -2019 6714 -1998 6730
rect -1946 6714 -1929 6730
rect -1873 6714 -1871 6748
rect -2240 6696 -2205 6714
rect -2171 6696 -2136 6714
rect -2102 6696 -2067 6714
rect -2033 6696 -1998 6714
rect -1964 6696 -1929 6714
rect -1895 6696 -1871 6714
rect -10447 6682 -1873 6696
rect -8092 6656 -8058 6682
rect -10604 6606 -10533 6622
rect -10570 6572 -10533 6606
rect -10604 6538 -10533 6572
rect -10570 6504 -10533 6538
rect -10604 6475 -10533 6504
rect -9748 6606 -9714 6622
rect -9748 6538 -9714 6572
rect -10604 6470 -10326 6475
rect -10570 6456 -10326 6470
rect -10570 6436 -10446 6456
rect -10604 6422 -10446 6436
rect -10412 6422 -10360 6456
rect -10604 6416 -10326 6422
rect -9748 6470 -9714 6504
rect -9748 6420 -9714 6436
rect -8092 6606 -8058 6622
rect -8092 6538 -8058 6572
rect -8092 6470 -8058 6498
rect -8092 6420 -8058 6436
rect -6436 6606 -6402 6622
rect -6436 6538 -6402 6572
rect -6436 6470 -6402 6504
rect -6436 6420 -6402 6436
rect -5580 6606 -5546 6622
rect -5580 6559 -5546 6572
rect -5580 6470 -5546 6504
rect -10559 6336 -10543 6370
rect -10509 6336 -10470 6370
rect -10413 6336 -10397 6370
rect -10333 6336 -10324 6370
rect -10290 6336 -10287 6370
rect -10253 6336 -10251 6370
rect -10217 6336 -10207 6370
rect -10144 6336 -10127 6370
rect -10071 6336 -10047 6370
rect -9997 6336 -9967 6370
rect -9923 6336 -9886 6370
rect -9849 6336 -9809 6370
rect -9771 6336 -9759 6370
rect -9703 6336 -9691 6370
rect -9653 6336 -9618 6370
rect -9584 6336 -9549 6370
rect -9511 6336 -9480 6370
rect -9438 6336 -9411 6370
rect -9365 6336 -9342 6370
rect -9292 6336 -9273 6370
rect -9219 6336 -9203 6370
rect -9146 6336 -9133 6370
rect -9073 6336 -9063 6370
rect -9000 6336 -8993 6370
rect -8927 6336 -8923 6370
rect -8889 6336 -8888 6370
rect -8854 6336 -8853 6370
rect -8819 6336 -8815 6370
rect -8749 6336 -8741 6370
rect -8679 6336 -8667 6370
rect -8609 6336 -8593 6370
rect -8539 6336 -8519 6370
rect -8469 6336 -8445 6370
rect -8399 6336 -8371 6370
rect -8329 6336 -8297 6370
rect -8259 6336 -8223 6370
rect -8189 6336 -8153 6370
rect -8115 6336 -8103 6370
rect -8047 6336 -8035 6370
rect -7997 6336 -7962 6370
rect -7927 6336 -7893 6370
rect -7853 6336 -7824 6370
rect -7779 6336 -7755 6370
rect -7705 6336 -7686 6370
rect -7631 6336 -7617 6370
rect -7557 6336 -7547 6370
rect -7483 6336 -7477 6370
rect -7409 6336 -7407 6370
rect -7373 6336 -7369 6370
rect -7303 6336 -7296 6370
rect -7233 6336 -7223 6370
rect -7163 6336 -7150 6370
rect -7093 6336 -7077 6370
rect -7023 6336 -7004 6370
rect -6953 6336 -6931 6370
rect -6883 6336 -6858 6370
rect -6813 6336 -6785 6370
rect -6743 6336 -6712 6370
rect -6673 6336 -6639 6370
rect -6603 6336 -6567 6370
rect -6532 6336 -6497 6370
rect -6459 6336 -6447 6370
rect -6391 6336 -6379 6370
rect -6341 6336 -6306 6370
rect -6268 6336 -6233 6370
rect -6195 6336 -6160 6370
rect -6122 6336 -6087 6370
rect -6049 6336 -6014 6370
rect -5976 6336 -5941 6370
rect -5903 6336 -5869 6370
rect -5829 6336 -5797 6370
rect -5755 6336 -5725 6370
rect -5681 6336 -5653 6370
rect -5607 6336 -5591 6370
rect -10294 6212 -10282 6246
rect -10244 6212 -10210 6246
rect -10176 6212 -10160 6246
rect -10339 6150 -10305 6162
rect -10339 6078 -10305 6112
rect -10339 6010 -10305 6044
rect -10339 5960 -10305 5972
rect -10163 6150 -10129 6162
rect -10163 6078 -10129 6112
rect -10163 6010 -10129 6044
rect -10163 5960 -10129 5972
<< viali >>
rect 6078 12672 6112 12706
rect 5823 12621 5857 12655
rect 5895 12621 5925 12655
rect 5925 12621 5929 12655
rect 6078 12600 6112 12634
rect 5776 12513 5810 12543
rect 5776 12509 5810 12513
rect 5776 12445 5810 12471
rect 5776 12437 5810 12445
rect 5958 12513 5986 12543
rect 5986 12513 5992 12543
rect 5958 12509 5992 12513
rect 5958 12445 5986 12471
rect 5986 12445 5992 12471
rect 5958 12437 5992 12445
rect 6314 12513 6344 12547
rect 6344 12513 6348 12547
rect 6314 12445 6344 12475
rect 6344 12445 6348 12475
rect 6314 12441 6348 12445
rect 5528 12303 5562 12337
rect 5528 12231 5562 12265
rect 5700 12143 5734 12177
rect 5700 12075 5734 12105
rect 5700 12071 5734 12075
rect 5856 12014 5860 12048
rect 5860 12014 5890 12048
rect 5986 12014 5996 12048
rect 5996 12014 6020 12048
rect 5700 11987 5734 11991
rect 5700 11957 5734 11987
rect 5700 11911 5734 11912
rect 5700 11878 5734 11911
rect 6248 11872 6282 11906
rect 5700 11800 5734 11833
rect 6248 11800 6282 11834
rect 5700 11799 5734 11800
rect 5700 11723 5734 11753
rect 5700 11719 5734 11723
rect 5856 11662 5860 11696
rect 5860 11662 5890 11696
rect 5986 11662 5996 11696
rect 5996 11662 6020 11696
rect 5700 11635 5734 11639
rect 5700 11605 5734 11635
rect 5700 11557 5734 11560
rect 5700 11526 5734 11557
rect 5700 11479 5734 11481
rect 5700 11447 5734 11479
rect 6163 11442 6197 11476
rect 5700 11367 5734 11401
rect 6163 11367 6197 11401
rect 5700 11289 5734 11321
rect 5700 11287 5734 11289
rect 5700 11211 5734 11241
rect 5700 11207 5734 11211
rect 5856 11150 5860 11184
rect 5860 11150 5890 11184
rect 5986 11150 5996 11184
rect 5996 11150 6020 11184
rect 5700 11123 5734 11127
rect 5700 11093 5734 11123
rect 5700 11045 5734 11048
rect 5700 11014 5734 11045
rect 5700 10967 5734 10969
rect 5700 10935 5734 10967
rect 6163 10930 6197 10964
rect 5700 10855 5734 10889
rect 6163 10855 6197 10889
rect 5700 10777 5734 10809
rect 5700 10775 5734 10777
rect 5700 10699 5734 10729
rect 5700 10695 5734 10699
rect 5856 10638 5860 10672
rect 5860 10638 5890 10672
rect 5986 10638 5996 10672
rect 5996 10638 6020 10672
rect 5700 10611 5734 10615
rect 5700 10581 5734 10611
rect 5700 10533 5734 10536
rect 5700 10502 5734 10533
rect 5700 10455 5734 10457
rect 5700 10423 5734 10455
rect 6078 10417 6112 10451
rect 5700 10343 5734 10377
rect 6078 10342 6112 10376
rect 5700 10265 5734 10297
rect 5700 10263 5734 10265
rect 5700 10187 5734 10217
rect 5700 10183 5734 10187
rect 5856 10126 5860 10160
rect 5860 10126 5890 10160
rect 5986 10126 5996 10160
rect 5996 10126 6020 10160
rect 5700 10099 5734 10103
rect 5700 10069 5734 10099
rect 5700 10021 5734 10024
rect 5700 9990 5734 10021
rect 5700 9943 5734 9945
rect 5700 9911 5734 9943
rect 6078 9905 6112 9939
rect 5700 9831 5734 9865
rect 6078 9830 6112 9864
rect 5700 9753 5734 9785
rect 5700 9751 5734 9753
rect 5700 9675 5734 9705
rect 5700 9671 5734 9675
rect 5856 9614 5860 9648
rect 5860 9614 5890 9648
rect 5986 9614 5996 9648
rect 5996 9614 6020 9648
rect 5772 9566 5806 9600
rect 5772 9494 5806 9528
rect 5913 9386 5947 9408
rect 5913 9374 5947 9386
rect 5913 9250 5947 9278
rect 6075 9420 6109 9423
rect 6075 9389 6089 9420
rect 6089 9389 6109 9420
rect 6075 9284 6109 9302
rect 6075 9268 6089 9284
rect 6089 9268 6109 9284
rect 5913 9244 5947 9250
rect 5969 9150 5974 9178
rect 5974 9150 6003 9178
rect 6043 9150 6050 9178
rect 6050 9150 6077 9178
rect 5969 9144 6003 9150
rect 6043 9144 6077 9150
rect 5606 9072 5640 9106
rect 6333 9072 6367 9106
rect 5606 9000 5640 9034
rect 6333 9000 6367 9034
rect 5778 8906 5812 8940
rect 6249 8883 6283 8917
rect 5778 8834 5812 8868
rect 6249 8810 6283 8844
rect -10534 7874 -10500 7908
rect -10462 7902 -10428 7908
rect -10462 7874 -10444 7902
rect -10444 7874 -10428 7902
rect -10382 7859 -10348 7893
rect -10382 7807 -10350 7808
rect -10350 7807 -10348 7808
rect -10382 7774 -10348 7807
rect -10382 7689 -10348 7723
rect -10382 7604 -10348 7638
rect -10382 7519 -10348 7553
rect -10262 7887 -10228 7893
rect -10262 7859 -10228 7887
rect -10262 7785 -10228 7808
rect -10262 7774 -10228 7785
rect -10262 7717 -10228 7723
rect -10262 7689 -10228 7717
rect -10262 7615 -10228 7638
rect -10262 7604 -10228 7615
rect -10262 7547 -10228 7553
rect -10262 7519 -10228 7547
rect -10086 7649 -10052 7670
rect -10086 7636 -10052 7649
rect -10086 7581 -10052 7589
rect -10086 7555 -10052 7581
rect -10086 7479 -10052 7509
rect -10086 7475 -10052 7479
rect -9910 7989 -9876 7993
rect -9910 7959 -9876 7989
rect -9910 7887 -9876 7911
rect -9687 7987 -9653 7996
rect -9687 7962 -9662 7987
rect -9662 7962 -9653 7987
rect -9687 7890 -9653 7924
rect -9568 7926 -9534 7930
rect -9568 7896 -9534 7926
rect -9910 7877 -9876 7887
rect -9910 7819 -9876 7829
rect -9910 7795 -9876 7819
rect -9910 7717 -9876 7746
rect -9910 7712 -9876 7717
rect -9910 7649 -9876 7663
rect -9910 7629 -9876 7649
rect -9910 7547 -9876 7580
rect -9568 7820 -9534 7849
rect -9568 7815 -9534 7820
rect -9568 7748 -9534 7768
rect -9568 7734 -9534 7748
rect -9568 7676 -9534 7687
rect -9568 7653 -9534 7676
rect -9568 7604 -9534 7606
rect -9568 7572 -9534 7604
rect -9910 7546 -9876 7547
rect -9910 7479 -9876 7497
rect -9910 7463 -9876 7479
rect -9687 7538 -9653 7572
rect -9687 7497 -9662 7500
rect -9662 7497 -9653 7500
rect -9687 7466 -9653 7497
rect -9568 7494 -9534 7525
rect -9568 7491 -9534 7494
rect -10490 7446 -10456 7455
rect -10490 7421 -10478 7446
rect -10478 7421 -10456 7446
rect -10490 7349 -10456 7383
rect -9568 7422 -9534 7444
rect -9568 7410 -9534 7422
rect -10029 7353 -9995 7365
rect -9957 7353 -9923 7365
rect -10219 7319 -10215 7353
rect -10215 7319 -10185 7353
rect -10147 7319 -10113 7353
rect -10029 7331 -10025 7353
rect -10025 7331 -9995 7353
rect -9957 7331 -9923 7353
rect -9568 7350 -9534 7363
rect -9568 7329 -9534 7350
rect -10447 6714 -10442 6748
rect -10442 6714 -10413 6748
rect -10375 6714 -10341 6748
rect -10303 6714 -10269 6748
rect -10231 6714 -10197 6748
rect -10159 6714 -10125 6748
rect -10087 6714 -10053 6748
rect -10015 6714 -9981 6748
rect -9943 6714 -9909 6748
rect -9871 6714 -9837 6748
rect -9799 6714 -9765 6748
rect -9727 6714 -9693 6748
rect -9655 6714 -9621 6748
rect -9583 6714 -9549 6748
rect -9511 6714 -9477 6748
rect -9439 6714 -9405 6748
rect -9367 6714 -9333 6748
rect -9295 6714 -9261 6748
rect -9223 6714 -9189 6748
rect -9151 6714 -9117 6748
rect -9079 6714 -9045 6748
rect -9007 6714 -8973 6748
rect -8935 6714 -8901 6748
rect -8863 6714 -8829 6748
rect -8791 6714 -8757 6748
rect -8719 6714 -8685 6748
rect -8647 6714 -8613 6748
rect -8575 6714 -8541 6748
rect -8503 6714 -8469 6748
rect -8431 6714 -8397 6748
rect -8359 6714 -8325 6748
rect -8287 6714 -8253 6748
rect -8215 6714 -8181 6748
rect -8143 6714 -8109 6748
rect -8071 6714 -8037 6748
rect -7999 6714 -7965 6748
rect -7927 6714 -7893 6748
rect -7855 6714 -7821 6748
rect -7783 6714 -7749 6748
rect -7711 6714 -7677 6748
rect -7639 6714 -7605 6748
rect -7567 6714 -7533 6748
rect -7495 6714 -7461 6748
rect -7423 6714 -7389 6748
rect -7351 6714 -7317 6748
rect -7279 6714 -7245 6748
rect -7207 6714 -7173 6748
rect -7135 6714 -7101 6748
rect -7063 6714 -7029 6748
rect -6991 6714 -6957 6748
rect -6919 6714 -6885 6748
rect -6847 6714 -6813 6748
rect -6775 6714 -6741 6748
rect -6703 6714 -6669 6748
rect -6631 6714 -6597 6748
rect -6559 6714 -6525 6748
rect -6487 6714 -6453 6748
rect -6415 6714 -6381 6748
rect -6343 6714 -6309 6748
rect -6271 6714 -6237 6748
rect -6199 6714 -6165 6748
rect -6127 6714 -6093 6748
rect -6055 6714 -6021 6748
rect -5983 6714 -5949 6748
rect -5911 6714 -5877 6748
rect -5839 6714 -5805 6748
rect -5767 6714 -5733 6748
rect -5695 6714 -5661 6748
rect -5623 6714 -5589 6748
rect -5551 6714 -5517 6748
rect -5479 6714 -5445 6748
rect -5407 6714 -5373 6748
rect -5335 6714 -5301 6748
rect -5263 6714 -5229 6748
rect -5191 6714 -5157 6748
rect -5119 6714 -5085 6748
rect -5046 6714 -5012 6748
rect -4973 6714 -4939 6748
rect -4900 6714 -4866 6748
rect -4827 6714 -4793 6748
rect -4754 6714 -4720 6748
rect -4681 6714 -4647 6748
rect -4608 6714 -4574 6748
rect -4535 6714 -4501 6748
rect -4462 6714 -4428 6748
rect -4389 6714 -4355 6748
rect -4316 6714 -4282 6748
rect -4243 6714 -4209 6748
rect -4170 6714 -4136 6748
rect -4097 6714 -4063 6748
rect -4024 6714 -3990 6748
rect -3951 6714 -3917 6748
rect -3878 6714 -3844 6748
rect -3805 6714 -3771 6748
rect -3732 6714 -3698 6748
rect -3659 6714 -3625 6748
rect -3586 6714 -3552 6748
rect -3513 6714 -3479 6748
rect -3440 6714 -3406 6748
rect -3367 6714 -3333 6748
rect -3294 6714 -3260 6748
rect -3221 6714 -3187 6748
rect -3148 6714 -3114 6748
rect -3075 6714 -3041 6748
rect -3002 6714 -2968 6748
rect -2929 6714 -2895 6748
rect -2856 6714 -2822 6748
rect -2783 6730 -2749 6748
rect -2710 6730 -2676 6748
rect -2637 6730 -2603 6748
rect -2564 6730 -2530 6748
rect -2491 6730 -2457 6748
rect -2418 6730 -2384 6748
rect -2345 6730 -2311 6748
rect -2272 6730 -2238 6748
rect -2199 6730 -2165 6748
rect -2126 6730 -2092 6748
rect -2053 6730 -2019 6748
rect -1980 6730 -1946 6748
rect -1907 6730 -1873 6748
rect -2783 6714 -2757 6730
rect -2757 6714 -2749 6730
rect -2710 6714 -2688 6730
rect -2688 6714 -2676 6730
rect -2637 6714 -2619 6730
rect -2619 6714 -2603 6730
rect -2564 6714 -2550 6730
rect -2550 6714 -2530 6730
rect -2491 6714 -2481 6730
rect -2481 6714 -2457 6730
rect -2418 6714 -2412 6730
rect -2412 6714 -2384 6730
rect -2345 6714 -2343 6730
rect -2343 6714 -2311 6730
rect -2272 6714 -2240 6730
rect -2240 6714 -2238 6730
rect -2199 6714 -2171 6730
rect -2171 6714 -2165 6730
rect -2126 6714 -2102 6730
rect -2102 6714 -2092 6730
rect -2053 6714 -2033 6730
rect -2033 6714 -2019 6730
rect -1980 6714 -1964 6730
rect -1964 6714 -1946 6730
rect -1907 6714 -1895 6730
rect -1895 6714 -1873 6730
rect -8092 6622 -8058 6656
rect -10446 6422 -10412 6456
rect -10360 6422 -10326 6456
rect -8092 6504 -8058 6532
rect -8092 6498 -8058 6504
rect -5580 6538 -5546 6559
rect -5580 6525 -5546 6538
rect -5580 6436 -5546 6453
rect -5580 6419 -5546 6436
rect -10447 6336 -10436 6370
rect -10436 6336 -10413 6370
rect -10367 6336 -10363 6370
rect -10363 6336 -10333 6370
rect -10287 6336 -10253 6370
rect -10207 6336 -10178 6370
rect -10178 6336 -10173 6370
rect -10127 6336 -10105 6370
rect -10105 6336 -10093 6370
rect -10047 6336 -10031 6370
rect -10031 6336 -10013 6370
rect -9967 6336 -9957 6370
rect -9957 6336 -9933 6370
rect -9886 6336 -9883 6370
rect -9883 6336 -9852 6370
rect -9805 6336 -9775 6370
rect -9775 6336 -9771 6370
rect -9691 6336 -9687 6370
rect -9687 6336 -9657 6370
rect -9618 6336 -9584 6370
rect -9545 6336 -9515 6370
rect -9515 6336 -9511 6370
rect -9472 6336 -9446 6370
rect -9446 6336 -9438 6370
rect -9399 6336 -9377 6370
rect -9377 6336 -9365 6370
rect -9326 6336 -9308 6370
rect -9308 6336 -9292 6370
rect -9253 6336 -9239 6370
rect -9239 6336 -9219 6370
rect -9180 6336 -9169 6370
rect -9169 6336 -9146 6370
rect -9107 6336 -9099 6370
rect -9099 6336 -9073 6370
rect -9034 6336 -9029 6370
rect -9029 6336 -9000 6370
rect -8961 6336 -8959 6370
rect -8959 6336 -8927 6370
rect -8888 6336 -8854 6370
rect -8815 6336 -8783 6370
rect -8783 6336 -8781 6370
rect -8741 6336 -8713 6370
rect -8713 6336 -8707 6370
rect -8667 6336 -8643 6370
rect -8643 6336 -8633 6370
rect -8593 6336 -8573 6370
rect -8573 6336 -8559 6370
rect -8519 6336 -8503 6370
rect -8503 6336 -8485 6370
rect -8445 6336 -8433 6370
rect -8433 6336 -8411 6370
rect -8371 6336 -8363 6370
rect -8363 6336 -8337 6370
rect -8297 6336 -8293 6370
rect -8293 6336 -8263 6370
rect -8223 6336 -8189 6370
rect -8149 6336 -8119 6370
rect -8119 6336 -8115 6370
rect -8035 6336 -8031 6370
rect -8031 6336 -8001 6370
rect -7961 6336 -7928 6370
rect -7928 6336 -7927 6370
rect -7887 6336 -7859 6370
rect -7859 6336 -7853 6370
rect -7813 6336 -7790 6370
rect -7790 6336 -7779 6370
rect -7739 6336 -7721 6370
rect -7721 6336 -7705 6370
rect -7665 6336 -7652 6370
rect -7652 6336 -7631 6370
rect -7591 6336 -7583 6370
rect -7583 6336 -7557 6370
rect -7517 6336 -7513 6370
rect -7513 6336 -7483 6370
rect -7443 6336 -7409 6370
rect -7369 6336 -7337 6370
rect -7337 6336 -7335 6370
rect -7296 6336 -7267 6370
rect -7267 6336 -7262 6370
rect -7223 6336 -7197 6370
rect -7197 6336 -7189 6370
rect -7150 6336 -7127 6370
rect -7127 6336 -7116 6370
rect -7077 6336 -7057 6370
rect -7057 6336 -7043 6370
rect -7004 6336 -6987 6370
rect -6987 6336 -6970 6370
rect -6931 6336 -6917 6370
rect -6917 6336 -6897 6370
rect -6858 6336 -6847 6370
rect -6847 6336 -6824 6370
rect -6785 6336 -6777 6370
rect -6777 6336 -6751 6370
rect -6712 6336 -6707 6370
rect -6707 6336 -6678 6370
rect -6639 6336 -6637 6370
rect -6637 6336 -6605 6370
rect -6566 6336 -6533 6370
rect -6533 6336 -6532 6370
rect -6493 6336 -6463 6370
rect -6463 6336 -6459 6370
rect -6379 6336 -6375 6370
rect -6375 6336 -6345 6370
rect -6306 6336 -6302 6370
rect -6302 6336 -6272 6370
rect -6233 6336 -6229 6370
rect -6229 6336 -6199 6370
rect -6160 6336 -6156 6370
rect -6156 6336 -6126 6370
rect -6087 6336 -6083 6370
rect -6083 6336 -6053 6370
rect -6014 6336 -6010 6370
rect -6010 6336 -5980 6370
rect -5941 6336 -5937 6370
rect -5937 6336 -5907 6370
rect -5869 6336 -5863 6370
rect -5863 6336 -5835 6370
rect -5797 6336 -5789 6370
rect -5789 6336 -5763 6370
rect -5725 6336 -5715 6370
rect -5715 6336 -5691 6370
rect -5653 6336 -5641 6370
rect -5641 6336 -5619 6370
rect -10282 6212 -10278 6246
rect -10278 6212 -10248 6246
rect -10210 6212 -10176 6246
rect -10339 6146 -10305 6150
rect -10339 6116 -10305 6146
rect -10339 6044 -10305 6078
rect -10339 5976 -10305 6006
rect -10339 5972 -10305 5976
rect -10163 6146 -10129 6150
rect -10163 6116 -10129 6146
rect -10163 6044 -10129 6078
rect -10163 5976 -10129 6006
rect -10163 5972 -10129 5976
<< metal1 >>
rect 5690 12782 6248 12812
tri 6248 12782 6278 12812 sw
rect 5690 12776 6278 12782
rect 5742 12772 6278 12776
tri 6278 12772 6288 12782 sw
rect 5742 12766 6288 12772
tri 5742 12741 5767 12766 nw
tri 6210 12741 6235 12766 ne
rect 6235 12741 6288 12766
tri 6235 12734 6242 12741 ne
rect 5690 12712 5742 12724
rect 6154 12720 6206 12726
rect 6072 12706 6118 12718
rect 6072 12672 6078 12706
rect 6112 12672 6118 12706
rect 5813 12661 5819 12664
rect 5690 12654 5742 12660
rect 5811 12615 5819 12661
rect 5813 12612 5819 12615
rect 5871 12612 5883 12664
rect 5935 12612 5941 12664
rect 6072 12634 6118 12672
rect 6072 12600 6078 12634
rect 6112 12600 6118 12634
rect 5606 12543 5816 12555
rect 5606 12509 5776 12543
rect 5810 12509 5816 12543
rect 5606 12471 5816 12509
rect 5606 12437 5776 12471
rect 5810 12437 5816 12471
rect 5606 12425 5816 12437
rect 5844 12543 6032 12557
rect 5844 12509 5958 12543
rect 5992 12509 6032 12543
rect 5844 12471 6032 12509
rect 5844 12437 5958 12471
rect 5992 12437 6032 12471
rect 5522 12337 5568 12349
rect 5522 12303 5528 12337
rect 5562 12303 5568 12337
rect 5522 12265 5568 12303
rect 5522 12231 5528 12265
rect 5562 12231 5568 12265
rect 5522 8153 5568 12231
rect 5606 12014 5652 12425
rect 5694 12187 5740 12189
rect 5690 12181 5742 12187
rect 5690 12117 5742 12129
rect 5690 12059 5742 12065
rect 5844 12048 6032 12437
tri 5652 12014 5676 12038 sw
rect 5844 12014 5856 12048
rect 5890 12014 5986 12048
rect 6020 12014 6032 12048
rect 5606 12003 5676 12014
tri 5676 12003 5687 12014 sw
rect 5606 11991 5740 12003
rect 5606 11957 5700 11991
rect 5734 11957 5740 11991
rect 5606 11912 5740 11957
rect 5606 11878 5700 11912
rect 5734 11878 5740 11912
rect 5606 11833 5740 11878
rect 5606 11799 5700 11833
rect 5734 11799 5740 11833
rect 5606 11753 5740 11799
rect 5606 11719 5700 11753
rect 5734 11719 5740 11753
rect 5606 11707 5740 11719
rect 5606 11696 5674 11707
tri 5674 11696 5685 11707 nw
rect 5844 11696 6032 12014
rect 5606 9231 5652 11696
tri 5652 11674 5674 11696 nw
rect 5844 11662 5856 11696
rect 5890 11662 5986 11696
rect 6020 11662 6032 11696
rect 5694 11639 5740 11651
rect 5694 11605 5700 11639
rect 5734 11605 5740 11639
rect 5694 11560 5740 11605
rect 5694 11526 5700 11560
rect 5734 11526 5740 11560
rect 5694 11481 5740 11526
rect 5694 11447 5700 11481
rect 5734 11447 5740 11481
rect 5694 11401 5740 11447
rect 5694 11367 5700 11401
rect 5734 11367 5740 11401
rect 5694 11321 5740 11367
rect 5694 11287 5700 11321
rect 5734 11287 5740 11321
rect 5694 11241 5740 11287
rect 5694 11207 5700 11241
rect 5734 11207 5740 11241
rect 5694 11202 5740 11207
tri 5740 11202 5812 11274 sw
rect 5694 11195 5812 11202
tri 5740 11184 5751 11195 ne
rect 5751 11184 5812 11195
tri 5751 11162 5773 11184 ne
rect 5694 11127 5740 11139
rect 5694 11093 5700 11127
rect 5734 11093 5740 11127
rect 5694 11048 5740 11093
rect 5694 11014 5700 11048
rect 5734 11014 5740 11048
rect 5694 10969 5740 11014
rect 5694 10935 5700 10969
rect 5734 10935 5740 10969
rect 5694 10889 5740 10935
rect 5694 10855 5700 10889
rect 5734 10855 5740 10889
rect 5694 10846 5740 10855
rect 5688 10840 5740 10846
rect 5688 10776 5700 10788
rect 5734 10776 5740 10788
rect 5688 10718 5700 10724
rect 5694 10695 5700 10718
rect 5734 10695 5740 10724
rect 5694 10683 5740 10695
rect 5688 10622 5740 10628
rect 5688 10558 5740 10570
rect 5688 10502 5700 10506
rect 5734 10502 5740 10506
rect 5688 10500 5740 10502
rect 5694 10457 5740 10500
rect 5694 10423 5700 10457
rect 5734 10423 5740 10457
rect 5694 10377 5740 10423
rect 5694 10343 5700 10377
rect 5734 10343 5740 10377
rect 5694 10297 5740 10343
rect 5694 10263 5700 10297
rect 5734 10263 5740 10297
rect 5694 10217 5740 10263
rect 5694 10183 5700 10217
rect 5734 10183 5740 10217
rect 5694 10171 5740 10183
rect 5694 10103 5740 10115
rect 5694 10069 5700 10103
rect 5734 10069 5740 10103
rect 5694 10024 5740 10069
rect 5694 9990 5700 10024
rect 5734 9990 5740 10024
rect 5694 9945 5740 9990
rect 5694 9911 5700 9945
rect 5734 9911 5740 9945
rect 5694 9865 5740 9911
rect 5694 9831 5700 9865
rect 5734 9831 5740 9865
rect 5694 9785 5740 9831
rect 5694 9751 5700 9785
rect 5734 9751 5740 9785
rect 5694 9705 5740 9751
rect 5694 9671 5700 9705
rect 5734 9671 5740 9705
tri 5686 9659 5694 9667 se
rect 5694 9659 5740 9671
rect 5686 9434 5732 9659
tri 5732 9651 5740 9659 nw
rect 5773 9612 5812 11184
rect 5766 9600 5812 9612
rect 5766 9566 5772 9600
rect 5806 9566 5812 9600
rect 5766 9528 5812 9566
rect 5766 9494 5772 9528
rect 5806 9494 5812 9528
rect 5766 9482 5812 9494
rect 5844 11184 6032 11662
rect 5844 11150 5856 11184
rect 5890 11150 5986 11184
rect 6020 11150 6032 11184
rect 5844 10672 6032 11150
rect 6072 10846 6118 12600
rect 6154 12656 6206 12668
rect 6154 12598 6206 12604
rect 6157 11476 6203 12598
rect 6242 12559 6288 12741
tri 6288 12559 6325 12596 sw
rect 6242 12547 6373 12559
rect 6242 12513 6314 12547
rect 6348 12513 6373 12547
rect 6242 12475 6373 12513
rect 6242 12441 6314 12475
rect 6348 12441 6373 12475
rect 6242 12429 6373 12441
rect 6243 11918 6289 11924
rect 6242 11906 6289 11918
rect 6242 11872 6248 11906
rect 6282 11872 6289 11906
rect 6242 11834 6289 11872
rect 6242 11800 6248 11834
rect 6282 11800 6289 11834
rect 6242 11788 6289 11800
rect 6157 11442 6163 11476
rect 6197 11442 6203 11476
rect 6157 11401 6203 11442
rect 6157 11367 6163 11401
rect 6197 11367 6203 11401
rect 6157 10964 6203 11367
rect 6157 10930 6163 10964
rect 6197 10930 6203 10964
rect 6157 10889 6203 10930
rect 6157 10855 6163 10889
rect 6197 10855 6203 10889
rect 6069 10840 6121 10846
rect 6069 10776 6121 10788
rect 6069 10718 6121 10724
rect 5844 10638 5856 10672
rect 5890 10638 5986 10672
rect 6020 10638 6032 10672
rect 5844 10160 6032 10638
rect 5844 10126 5856 10160
rect 5890 10126 5986 10160
rect 6020 10126 6032 10160
rect 5844 10032 6032 10126
rect 5844 9980 5847 10032
rect 5899 9980 5911 10032
rect 5963 9980 5975 10032
rect 6027 9980 6032 10032
rect 5844 9950 6032 9980
rect 5844 9898 5847 9950
rect 5899 9898 5911 9950
rect 5963 9898 5975 9950
rect 6027 9898 6032 9950
rect 5844 9868 6032 9898
rect 5844 9816 5847 9868
rect 5899 9816 5911 9868
rect 5963 9816 5975 9868
rect 6027 9816 6032 9868
rect 5844 9785 6032 9816
rect 5844 9733 5847 9785
rect 5899 9733 5911 9785
rect 5963 9733 5975 9785
rect 6027 9733 6032 9785
rect 5844 9648 6032 9733
rect 5844 9614 5856 9648
rect 5890 9614 5986 9648
rect 6020 9614 6032 9648
rect 6072 10451 6118 10718
rect 6157 10628 6203 10855
rect 6154 10622 6206 10628
rect 6154 10558 6206 10570
rect 6154 10500 6206 10506
rect 6072 10417 6078 10451
rect 6112 10417 6118 10451
rect 6072 10376 6118 10417
rect 6072 10342 6078 10376
rect 6112 10342 6118 10376
rect 6072 9939 6118 10342
rect 6072 9905 6078 9939
rect 6112 9905 6118 9939
rect 6072 9864 6118 9905
rect 6072 9830 6078 9864
rect 6112 9830 6118 9864
rect 6072 9621 6118 9830
rect 5844 9526 6032 9614
rect 5844 9493 5999 9526
tri 5999 9493 6032 9526 nw
rect 6069 9615 6121 9621
rect 6069 9551 6121 9563
rect 6069 9493 6121 9499
tri 5732 9434 5756 9458 sw
rect 5686 9428 5756 9434
rect 5686 9376 5704 9428
rect 5686 9364 5756 9376
rect 5686 9312 5704 9364
rect 5686 9306 5756 9312
rect 5844 9408 5964 9493
tri 5964 9458 5999 9493 nw
rect 6157 9445 6203 10500
rect 6157 9439 6209 9445
rect 6069 9434 6115 9435
rect 5844 9374 5913 9408
rect 5947 9374 5964 9408
rect 5844 9278 5964 9374
rect 6066 9428 6118 9434
rect 6066 9364 6118 9376
rect 6157 9375 6209 9387
rect 6157 9317 6209 9323
rect 6066 9306 6118 9312
tri 6118 9306 6123 9311 sw
rect 5844 9244 5913 9278
rect 5947 9244 5964 9278
rect 6069 9302 6123 9306
rect 6069 9268 6075 9302
rect 6109 9268 6123 9302
rect 6069 9256 6123 9268
tri 6123 9256 6173 9306 sw
tri 5652 9231 5657 9236 sw
rect 5844 9231 5964 9244
tri 6080 9241 6095 9256 ne
rect 6095 9241 6173 9256
tri 6173 9241 6188 9256 sw
tri 6095 9231 6105 9241 ne
rect 6105 9231 6188 9241
rect 5606 9222 5657 9231
tri 5657 9222 5666 9231 sw
tri 6105 9222 6114 9231 ne
rect 6114 9222 6188 9231
rect 5606 9209 5666 9222
tri 5606 9207 5608 9209 ne
rect 5608 9207 5666 9209
tri 5666 9207 5681 9222 sw
tri 6114 9207 6129 9222 ne
rect 6129 9207 6188 9222
tri 5608 9178 5637 9207 ne
rect 5637 9200 5681 9207
tri 5681 9200 5688 9207 sw
tri 6129 9200 6136 9207 ne
rect 5637 9184 5688 9200
tri 5688 9184 5704 9200 sw
rect 5637 9178 5704 9184
tri 5704 9178 5710 9184 sw
rect 5957 9178 6089 9184
tri 5637 9163 5652 9178 ne
rect 5652 9163 5710 9178
tri 5652 9144 5671 9163 ne
rect 5671 9144 5710 9163
tri 5710 9144 5744 9178 sw
rect 5957 9144 5969 9178
rect 6003 9144 6043 9178
rect 6077 9144 6089 9178
tri 5671 9134 5681 9144 ne
rect 5681 9138 5744 9144
tri 5744 9138 5750 9144 sw
rect 5957 9138 6089 9144
rect 5681 9134 5750 9138
tri 5750 9134 5754 9138 sw
tri 5681 9119 5696 9134 ne
rect 5696 9119 5754 9134
tri 5754 9119 5769 9134 sw
rect -10546 8061 -10457 8113
rect -10405 8061 -10391 8113
rect -10339 8061 -10333 8113
rect -9494 8107 -9442 8113
rect -10546 8008 -10410 8061
tri -10410 8008 -10357 8061 nw
rect 5424 8101 5430 8153
rect 5482 8101 5494 8153
rect 5546 8117 5568 8153
rect 5546 8113 5564 8117
tri 5564 8113 5568 8117 nw
rect 5600 9106 5652 9119
tri 5696 9106 5709 9119 ne
rect 5709 9106 5769 9119
tri 5769 9106 5782 9119 sw
rect 5600 9072 5606 9106
rect 5640 9072 5652 9106
tri 5709 9072 5743 9106 ne
rect 5743 9088 5782 9106
tri 5782 9088 5800 9106 sw
rect 5743 9072 5800 9088
tri 5800 9072 5816 9088 sw
rect 5931 9082 5983 9088
rect 5600 9034 5652 9072
tri 5743 9061 5754 9072 ne
rect 5754 9061 5816 9072
tri 5816 9061 5827 9072 sw
tri 5754 9034 5781 9061 ne
rect 5781 9034 5827 9061
tri 5827 9034 5854 9061 sw
rect 5600 9000 5606 9034
rect 5640 9000 5652 9034
tri 5781 9011 5804 9034 ne
rect 5804 9011 5854 9034
tri 5854 9011 5877 9034 sw
rect 5931 9018 5983 9030
rect 5546 8107 5558 8113
tri 5558 8107 5564 8113 nw
rect 5546 8101 5552 8107
tri 5552 8101 5558 8107 nw
rect 5600 8069 5652 9000
rect -9494 8041 -9442 8055
rect -10546 7908 -10416 8008
tri -10416 8002 -10410 8008 nw
rect -10546 7874 -10534 7908
rect -10500 7874 -10462 7908
rect -10428 7874 -10416 7908
rect -9916 7993 -9870 8005
rect -9916 7959 -9910 7993
rect -9876 7959 -9870 7993
rect -9916 7911 -9870 7959
rect -10546 7868 -10416 7874
rect -10388 7893 -10222 7905
rect -10388 7859 -10382 7893
rect -10348 7859 -10262 7893
rect -10228 7859 -10222 7893
rect -9916 7877 -9910 7911
rect -9876 7877 -9870 7911
rect -9696 8002 -9644 8008
rect 5508 8017 5514 8069
rect 5566 8017 5578 8069
rect 5630 8032 5652 8069
rect 5630 8017 5637 8032
tri 5637 8017 5652 8032 nw
rect 5684 9005 5736 9011
tri 5804 9000 5815 9011 ne
rect 5815 9000 5877 9011
tri 5877 9000 5888 9011 sw
tri 5815 8988 5827 9000 ne
rect 5827 8988 5888 9000
tri 5888 8988 5900 9000 sw
tri 5827 8967 5848 8988 ne
rect 5848 8979 5900 8988
rect 5684 8941 5736 8953
rect -9494 7983 -9442 7989
rect 5684 7985 5736 8889
tri -9494 7980 -9491 7983 ne
rect -9491 7980 -9445 7983
tri -9445 7980 -9442 7983 nw
tri -9491 7977 -9488 7980 ne
rect -9696 7936 -9644 7950
rect -9696 7878 -9644 7884
rect -9574 7930 -9522 7942
rect -9574 7896 -9568 7930
rect -9534 7896 -9522 7930
rect -10388 7849 -10222 7859
tri -10010 7854 -9999 7865 se
rect -9999 7859 -9947 7865
tri -10222 7849 -10217 7854 sw
tri -10015 7849 -10010 7854 se
rect -10010 7849 -9999 7854
rect -10388 7829 -10217 7849
tri -10217 7829 -10197 7849 sw
tri -10035 7829 -10015 7849 se
rect -10015 7829 -9999 7849
rect -10388 7825 -10197 7829
tri -10197 7825 -10193 7829 sw
tri -10039 7825 -10035 7829 se
rect -10035 7825 -9999 7829
rect -10388 7808 -9999 7825
rect -10388 7774 -10382 7808
rect -10348 7774 -10262 7808
rect -10228 7807 -9999 7808
rect -10228 7793 -9947 7807
rect -10228 7774 -9999 7793
rect -10388 7741 -9999 7774
rect -9916 7829 -9870 7877
rect -9916 7795 -9910 7829
rect -9876 7795 -9870 7829
rect -9916 7746 -9870 7795
rect -9916 7744 -9910 7746
rect -10388 7735 -9947 7741
rect -9919 7738 -9910 7744
rect -9876 7744 -9870 7746
rect -9574 7849 -9522 7896
rect -9574 7815 -9568 7849
rect -9534 7815 -9522 7849
rect -9574 7768 -9522 7815
rect -9876 7738 -9867 7744
rect -10388 7723 -10222 7735
rect -10388 7689 -10382 7723
rect -10348 7689 -10262 7723
rect -10228 7689 -10222 7723
rect -10388 7638 -10222 7689
rect -10388 7604 -10382 7638
rect -10348 7604 -10262 7638
rect -10228 7604 -10222 7638
rect -10092 7670 -10046 7682
rect -10092 7637 -10086 7670
rect -10388 7553 -10222 7604
rect -10388 7519 -10382 7553
rect -10348 7519 -10262 7553
rect -10228 7519 -10222 7553
rect -10388 7507 -10222 7519
rect -10095 7636 -10086 7637
rect -10052 7637 -10046 7670
rect -9919 7672 -9867 7686
rect -10052 7636 -10043 7637
rect -10095 7631 -10043 7636
rect -9919 7614 -9867 7620
rect -9574 7738 -9568 7768
rect -9534 7738 -9522 7768
rect -9574 7672 -9568 7686
rect -9534 7672 -9522 7686
rect -10095 7567 -10086 7579
rect -10052 7567 -10043 7579
tri -10097 7509 -10095 7511 se
rect -10095 7509 -10043 7515
rect -9916 7580 -9870 7614
rect -9574 7606 -9522 7620
rect -9916 7546 -9910 7580
rect -9876 7546 -9870 7580
tri -10099 7507 -10097 7509 se
rect -10097 7507 -10086 7509
tri -10131 7475 -10099 7507 se
rect -10099 7475 -10086 7507
rect -10052 7475 -10046 7509
tri -10139 7467 -10131 7475 se
rect -10131 7467 -10046 7475
rect -10505 7461 -10046 7467
rect -10453 7419 -10046 7461
rect -9916 7497 -9870 7546
rect -9916 7463 -9910 7497
rect -9876 7463 -9870 7497
rect -9916 7451 -9870 7463
rect -9696 7578 -9644 7584
rect -9696 7512 -9644 7526
rect -9696 7454 -9644 7460
rect -9574 7572 -9568 7606
rect -9534 7572 -9522 7606
rect -9574 7525 -9522 7572
rect -9574 7491 -9568 7525
rect -9534 7491 -9522 7525
rect -9574 7451 -9522 7491
rect -10453 7410 -10055 7419
tri -10055 7410 -10046 7419 nw
rect -10453 7409 -10068 7410
rect -10505 7397 -10068 7409
tri -10068 7397 -10055 7410 nw
rect -10453 7365 -10422 7397
tri -10422 7365 -10390 7397 nw
rect -9574 7385 -9522 7399
rect -10453 7353 -10434 7365
tri -10434 7353 -10422 7365 nw
rect -10453 7345 -10450 7353
rect -10505 7337 -10450 7345
tri -10450 7337 -10434 7353 nw
rect -10231 7307 -10225 7359
rect -10173 7307 -10161 7359
rect -10109 7307 -10101 7359
tri -10101 7307 -10085 7323 sw
rect -10041 7319 -10035 7371
rect -9983 7319 -9969 7371
rect -9917 7319 -9911 7371
rect -9686 7332 -9634 7338
tri -9691 7319 -9686 7324 se
tri -9703 7307 -9691 7319 se
rect -9691 7307 -9686 7319
rect -10231 7301 -10085 7307
tri -10085 7301 -10079 7307 sw
tri -9709 7301 -9703 7307 se
rect -9703 7301 -9686 7307
rect -10231 7291 -10079 7301
tri -10079 7291 -10069 7301 sw
tri -9719 7291 -9709 7301 se
rect -9709 7291 -9686 7301
rect -10231 7280 -9686 7291
rect -9574 7329 -9568 7333
rect -9534 7329 -9522 7333
rect -9574 7317 -9522 7329
rect -10231 7266 -9634 7280
rect -10231 7254 -9686 7266
tri -9718 7222 -9686 7254 ne
rect -9686 7208 -9634 7214
tri -9491 7174 -9488 7177 se
rect -9488 7174 -9445 7980
rect 5592 7933 5598 7985
rect 5650 7933 5662 7985
rect 5714 7949 5736 7985
rect 5714 7933 5720 7949
tri 5720 7933 5736 7949 nw
rect 5767 8940 5819 8955
rect 5767 8906 5778 8940
rect 5812 8906 5819 8940
rect 5767 8868 5819 8906
rect 5767 8834 5778 8868
rect 5812 8834 5819 8868
rect 5767 7901 5819 8834
rect 5675 7849 5681 7901
rect 5733 7849 5745 7901
rect 5797 7865 5819 7901
rect 5797 7849 5803 7865
tri 5803 7849 5819 7865 nw
rect 5848 8915 5900 8927
rect 5848 7817 5900 8863
rect 5755 7765 5761 7817
rect 5813 7765 5825 7817
rect 5877 7780 5900 7817
rect 5877 7765 5885 7780
tri 5885 7765 5900 7780 nw
rect 5931 7733 5983 8966
rect 5855 7681 5861 7733
rect 5913 7681 5925 7733
rect 5977 7681 5983 7733
rect 6025 8947 6077 9138
rect 6025 8883 6077 8895
rect 6025 7649 6077 8831
rect 5949 7597 5955 7649
rect 6007 7597 6019 7649
rect 6071 7597 6077 7649
rect 6136 7565 6188 9207
rect 6243 8917 6289 11788
rect 6327 9106 6373 12429
rect 6327 9072 6333 9106
rect 6367 9072 6373 9106
rect 6327 9034 6373 9072
rect 6327 9000 6333 9034
rect 6367 9000 6373 9034
rect 6327 8988 6373 9000
rect 6243 8883 6249 8917
rect 6283 8883 6289 8917
rect 6243 8844 6289 8883
rect 6243 8810 6249 8844
rect 6283 8810 6289 8844
rect 6243 8798 6289 8810
rect 6060 7513 6066 7565
rect 6118 7513 6130 7565
rect 6182 7513 6188 7565
tri -9445 7174 -9442 7177 sw
tri -9494 7171 -9491 7174 se
rect -9491 7171 -9442 7174
rect -9494 7165 -9442 7171
rect -9494 7099 -9442 7113
rect -9494 7041 -9442 7047
rect -10459 6748 -1861 6786
rect -10407 6714 -10375 6748
rect -10341 6714 -10303 6748
rect -10269 6714 -10231 6748
rect -10197 6714 -10159 6748
rect -10125 6714 -10087 6748
rect -10053 6714 -10015 6748
rect -9981 6714 -9943 6748
rect -9909 6714 -9871 6748
rect -9837 6714 -9799 6748
rect -9765 6714 -9727 6748
rect -9693 6714 -9655 6748
rect -9621 6714 -9583 6748
rect -9549 6714 -9511 6748
rect -9477 6714 -9439 6748
rect -9405 6714 -9367 6748
rect -9333 6714 -9295 6748
rect -9261 6714 -9223 6748
rect -9189 6714 -9151 6748
rect -9117 6714 -9079 6748
rect -9045 6714 -9007 6748
rect -8973 6714 -8935 6748
rect -8901 6714 -8863 6748
rect -8829 6714 -8791 6748
rect -8757 6714 -8719 6748
rect -8685 6714 -8647 6748
rect -8613 6714 -8575 6748
rect -8541 6714 -8503 6748
rect -8469 6714 -8431 6748
rect -8397 6714 -8359 6748
rect -8325 6714 -8287 6748
rect -8253 6714 -8215 6748
rect -8181 6714 -8143 6748
rect -8109 6714 -8071 6748
rect -8037 6714 -7999 6748
rect -7965 6714 -7927 6748
rect -7893 6714 -7855 6748
rect -7821 6714 -7783 6748
rect -7749 6714 -7711 6748
rect -7677 6714 -7639 6748
rect -7605 6714 -7567 6748
rect -7533 6714 -7495 6748
rect -7461 6714 -7423 6748
rect -7389 6714 -7351 6748
rect -7317 6714 -7279 6748
rect -7245 6714 -7207 6748
rect -7173 6714 -7135 6748
rect -7101 6714 -7063 6748
rect -7029 6714 -6991 6748
rect -6957 6714 -6919 6748
rect -6885 6714 -6847 6748
rect -6813 6714 -6775 6748
rect -6741 6714 -6703 6748
rect -6669 6714 -6631 6748
rect -6597 6714 -6559 6748
rect -6525 6714 -6487 6748
rect -6453 6714 -6415 6748
rect -6381 6714 -6343 6748
rect -6309 6714 -6271 6748
rect -6237 6714 -6199 6748
rect -6165 6714 -6127 6748
rect -6093 6714 -6055 6748
rect -6021 6714 -5983 6748
rect -5949 6714 -5911 6748
rect -5877 6714 -5839 6748
rect -5805 6714 -5767 6748
rect -5733 6714 -5695 6748
rect -5661 6714 -5623 6748
rect -5589 6714 -5551 6748
rect -5517 6714 -5479 6748
rect -5445 6714 -5407 6748
rect -5373 6714 -5335 6748
rect -5301 6714 -5263 6748
rect -5229 6714 -5191 6748
rect -5157 6714 -5119 6748
rect -5085 6714 -5046 6748
rect -5012 6714 -4973 6748
rect -4939 6714 -4900 6748
rect -4866 6714 -4827 6748
rect -4793 6714 -4754 6748
rect -4720 6714 -4681 6748
rect -4647 6714 -4608 6748
rect -4574 6714 -4535 6748
rect -4501 6714 -4462 6748
rect -4428 6714 -4389 6748
rect -4355 6714 -4316 6748
rect -4282 6714 -4243 6748
rect -4209 6714 -4170 6748
rect -4136 6714 -4097 6748
rect -4063 6714 -4024 6748
rect -3990 6714 -3951 6748
rect -3917 6714 -3878 6748
rect -3844 6714 -3805 6748
rect -3771 6714 -3732 6748
rect -3698 6714 -3659 6748
rect -3625 6714 -3586 6748
rect -3552 6714 -3513 6748
rect -3479 6714 -3440 6748
rect -3406 6714 -3367 6748
rect -3333 6714 -3294 6748
rect -3260 6714 -3221 6748
rect -3187 6714 -3148 6748
rect -3114 6714 -3075 6748
rect -3041 6714 -3002 6748
rect -2968 6714 -2929 6748
rect -2895 6714 -2856 6748
rect -2822 6714 -2783 6748
rect -2749 6714 -2710 6748
rect -2676 6714 -2637 6748
rect -2603 6714 -2564 6748
rect -2530 6714 -2491 6748
rect -2457 6714 -2418 6748
rect -2384 6714 -2345 6748
rect -2311 6714 -2272 6748
rect -2238 6714 -2199 6748
rect -2165 6714 -2126 6748
rect -2092 6714 -2053 6748
rect -2019 6714 -1980 6748
rect -1946 6714 -1907 6748
rect -1873 6714 -1861 6748
rect -10407 6696 -1861 6714
rect -10459 6679 -1861 6696
rect -10407 6676 -1861 6679
rect -10407 6656 -1886 6676
rect -10407 6627 -8092 6656
rect -10459 6622 -8092 6627
rect -8058 6622 -1886 6656
rect -10459 6610 -1886 6622
rect -10407 6599 -1886 6610
rect -10407 6571 -5694 6599
tri -5694 6571 -5666 6599 nw
tri -3765 6584 -3750 6599 ne
rect -3750 6584 -1886 6599
rect -10407 6559 -5706 6571
tri -5706 6559 -5694 6571 nw
rect -5586 6559 -5540 6571
rect -10407 6558 -5712 6559
rect -10459 6553 -5712 6558
tri -5712 6553 -5706 6559 nw
rect -10459 6552 -10407 6553
rect -8098 6532 -8052 6553
rect -8098 6498 -8092 6532
rect -8058 6498 -8052 6532
rect -8098 6486 -8052 6498
rect -5586 6525 -5580 6559
rect -5546 6554 -5540 6559
tri -5540 6554 -5523 6571 sw
rect -5546 6525 -5431 6554
tri -5590 6486 -5586 6490 se
rect -5586 6486 -5431 6525
tri -5608 6468 -5590 6486 se
rect -5590 6468 -5431 6486
tri -9986 6462 -9980 6468 se
rect -9980 6462 -9971 6468
rect -10459 6458 -10314 6462
tri -10314 6458 -10310 6462 sw
tri -9990 6458 -9986 6462 se
rect -9986 6458 -9971 6462
rect -10459 6456 -9971 6458
rect -10459 6422 -10446 6456
rect -10412 6422 -10360 6456
rect -10326 6422 -9971 6456
rect -10459 6416 -9971 6422
rect -9919 6416 -9898 6468
rect -9846 6462 -9810 6468
tri -9810 6462 -9804 6468 sw
tri -5614 6462 -5608 6468 se
rect -5608 6462 -5431 6468
rect -9846 6458 -9804 6462
tri -9804 6458 -9800 6462 sw
tri -5618 6458 -5614 6462 se
rect -5614 6458 -5431 6462
rect -9846 6416 -9233 6458
tri -9823 6407 -9814 6416 ne
rect -9814 6407 -9233 6416
tri -9814 6406 -9813 6407 ne
rect -9813 6406 -9233 6407
rect -9181 6406 -9160 6458
rect -9108 6406 -9102 6458
tri -8118 6453 -8113 6458 se
rect -8113 6453 -5431 6458
tri -8152 6419 -8118 6453 se
rect -8118 6419 -5580 6453
rect -5546 6419 -5431 6453
tri -8164 6407 -8152 6419 se
rect -8152 6407 -5431 6419
tri -8165 6406 -8164 6407 se
rect -8164 6406 -5431 6407
tri -8189 6382 -8165 6406 se
rect -8165 6382 -8097 6406
tri -8097 6382 -8073 6406 nw
tri -5586 6382 -5562 6406 ne
rect -5562 6382 -5431 6406
rect -9977 6376 -9971 6382
rect -10459 6370 -9971 6376
rect -10459 6336 -10447 6370
rect -10413 6336 -10367 6370
rect -10333 6336 -10287 6370
rect -10253 6336 -10207 6370
rect -10173 6336 -10127 6370
rect -10093 6336 -10047 6370
rect -10013 6336 -9971 6370
rect -10459 6330 -9971 6336
rect -9919 6330 -9898 6382
rect -9846 6376 -9840 6382
tri -8195 6376 -8189 6382 se
rect -8189 6376 -8103 6382
tri -8103 6376 -8097 6382 nw
tri -5562 6379 -5559 6382 ne
rect -9846 6370 -9759 6376
rect -9846 6336 -9805 6370
rect -9771 6336 -9759 6370
rect -9846 6330 -9759 6336
rect -9703 6370 -9664 6376
rect -9612 6370 -9591 6376
rect -9539 6370 -8103 6376
rect -9703 6336 -9691 6370
rect -9511 6336 -9472 6370
rect -9438 6336 -9399 6370
rect -9365 6336 -9326 6370
rect -9292 6336 -9253 6370
rect -9219 6336 -9180 6370
rect -9146 6336 -9107 6370
rect -9073 6336 -9034 6370
rect -9000 6336 -8961 6370
rect -8927 6336 -8888 6370
rect -8854 6336 -8815 6370
rect -8781 6336 -8741 6370
rect -8707 6336 -8667 6370
rect -8633 6336 -8593 6370
rect -8559 6336 -8519 6370
rect -8485 6336 -8445 6370
rect -8411 6336 -8371 6370
rect -8337 6336 -8297 6370
rect -8263 6336 -8223 6370
rect -8189 6336 -8149 6370
rect -8115 6336 -8103 6370
rect -9703 6330 -9664 6336
rect -9670 6324 -9664 6330
rect -9612 6324 -9591 6336
rect -9539 6330 -8103 6336
rect -9539 6324 -9533 6330
rect -8047 6324 -8041 6376
rect -7989 6324 -7968 6376
rect -7916 6370 -6447 6376
rect -7916 6336 -7887 6370
rect -7853 6336 -7813 6370
rect -7779 6336 -7739 6370
rect -7705 6336 -7665 6370
rect -7631 6336 -7591 6370
rect -7557 6336 -7517 6370
rect -7483 6336 -7443 6370
rect -7409 6336 -7369 6370
rect -7335 6336 -7296 6370
rect -7262 6336 -7223 6370
rect -7189 6336 -7150 6370
rect -7116 6336 -7077 6370
rect -7043 6336 -7004 6370
rect -6970 6336 -6931 6370
rect -6897 6336 -6858 6370
rect -6824 6336 -6785 6370
rect -6751 6336 -6712 6370
rect -6678 6336 -6639 6370
rect -6605 6336 -6566 6370
rect -6532 6336 -6493 6370
rect -6459 6336 -6447 6370
rect -7916 6330 -6447 6336
rect -6391 6370 -6186 6376
rect -6134 6370 -6113 6376
rect -6061 6370 -5607 6376
rect -6391 6336 -6379 6370
rect -6345 6336 -6306 6370
rect -6272 6336 -6233 6370
rect -6199 6336 -6186 6370
rect -6126 6336 -6113 6370
rect -6053 6336 -6014 6370
rect -5980 6336 -5941 6370
rect -5907 6336 -5869 6370
rect -5835 6336 -5797 6370
rect -5763 6336 -5725 6370
rect -5691 6336 -5653 6370
rect -5619 6336 -5607 6370
rect -6391 6330 -6186 6336
rect -7916 6324 -7910 6330
tri -6397 6324 -6391 6330 se
rect -6391 6324 -6343 6330
tri -6425 6296 -6397 6324 se
rect -6397 6296 -6343 6324
tri -6343 6296 -6309 6330 nw
rect -6192 6324 -6186 6330
rect -6134 6324 -6113 6336
rect -6061 6330 -5607 6336
rect -5559 6348 -5431 6382
rect -6061 6324 -6055 6330
rect -5559 6296 -5553 6348
rect -5501 6296 -5489 6348
rect -5437 6296 -5431 6348
tri -10098 6270 -10072 6296 se
rect -10072 6270 -6369 6296
tri -6369 6270 -6343 6296 nw
tri -3753 6270 -3736 6287 se
rect -3736 6270 -3730 6287
rect -10294 6256 -6383 6270
tri -6383 6256 -6369 6270 nw
tri -3767 6256 -3753 6270 se
rect -3753 6256 -3730 6270
rect -10294 6246 -10067 6256
rect -10294 6212 -10282 6246
rect -10248 6212 -10210 6246
rect -10176 6216 -10067 6246
tri -10067 6216 -10027 6256 nw
tri -3800 6223 -3767 6256 se
rect -3767 6235 -3730 6256
rect -3678 6235 -3666 6287
rect -3614 6235 -3608 6287
rect -3767 6223 -3736 6235
rect -10176 6215 -10068 6216
tri -10068 6215 -10067 6216 nw
rect -10176 6212 -10077 6215
rect -10294 6206 -10077 6212
tri -10077 6206 -10068 6215 nw
tri -11144 6192 -11141 6195 ne
rect -9239 6171 -9233 6223
rect -9181 6171 -9160 6223
rect -9108 6216 -9102 6223
tri -9102 6216 -9095 6223 sw
tri -8054 6216 -8047 6223 se
rect -8047 6216 -8041 6223
rect -9108 6215 -9095 6216
tri -9095 6215 -9094 6216 sw
tri -8055 6215 -8054 6216 se
rect -8054 6215 -8041 6216
rect -9108 6206 -9094 6215
tri -9094 6206 -9085 6215 sw
tri -8064 6206 -8055 6215 se
rect -8055 6206 -8041 6215
rect -9108 6203 -9085 6206
tri -9085 6203 -9082 6206 sw
tri -8067 6203 -8064 6206 se
rect -8064 6203 -8041 6206
rect -9108 6171 -8041 6203
rect -7989 6171 -7968 6223
rect -7916 6216 -7910 6223
tri -7910 6216 -7903 6223 sw
tri -3807 6216 -3800 6223 se
rect -3800 6216 -3736 6223
rect -7916 6215 -7903 6216
tri -7903 6215 -7902 6216 sw
tri -3808 6215 -3807 6216 se
rect -3807 6215 -3736 6216
tri -3736 6215 -3716 6235 nw
rect -7916 6203 -3748 6215
tri -3748 6203 -3736 6215 nw
rect -7916 6195 -3756 6203
tri -3756 6195 -3748 6203 nw
rect -7916 6192 -3759 6195
tri -3759 6192 -3756 6195 nw
rect -7916 6171 -3780 6192
tri -3780 6171 -3759 6192 nw
rect -10459 6156 -10299 6162
rect -10407 6150 -10299 6156
rect -10407 6116 -10339 6150
rect -10305 6116 -10299 6150
rect -10407 6104 -10299 6116
rect -10459 6087 -10299 6104
rect -10407 6078 -10299 6087
rect -10407 6044 -10339 6078
rect -10305 6044 -10299 6078
rect -10407 6035 -10299 6044
rect -10459 6018 -10299 6035
rect -10407 6006 -10299 6018
rect -10407 5972 -10339 6006
rect -10305 5972 -10299 6006
rect -10407 5966 -10299 5972
rect -10459 5960 -10299 5966
rect -10169 6150 -10123 6162
rect -10169 6116 -10163 6150
rect -10129 6116 -10123 6150
rect -10169 6078 -10123 6116
rect -10169 6044 -10163 6078
rect -10129 6060 -10123 6078
rect -9977 6131 -9925 6137
rect -9806 6110 -9800 6162
rect -9748 6110 -9727 6162
rect -9675 6142 -9669 6162
tri -9669 6142 -9649 6162 sw
rect -9675 6137 -5416 6142
tri -5416 6137 -5411 6142 sw
rect -9675 6110 -5411 6137
tri -5456 6103 -5449 6110 ne
rect -5449 6103 -5411 6110
tri -5411 6103 -5377 6137 sw
rect -9977 6066 -9925 6079
tri -5449 6070 -5416 6103 ne
rect -5416 6070 -5365 6103
rect -10129 6044 -9977 6060
rect -10169 6014 -9977 6044
tri -5416 6060 -5406 6070 ne
rect -5406 6060 -5365 6070
rect -9925 6014 -6886 6060
rect -10169 6008 -6886 6014
rect -6834 6008 -6817 6060
rect -6765 6008 -6748 6060
rect -6696 6008 -6690 6060
tri -5406 6051 -5397 6060 ne
rect -5397 6051 -5365 6060
rect -5313 6051 -5292 6103
rect -5240 6051 -5219 6103
rect -5167 6051 -5146 6103
rect -5094 6051 -5088 6103
rect -10169 6006 -10123 6008
rect -10169 5972 -10163 6006
rect -10129 5972 -10123 6006
rect -10169 5960 -10123 5972
<< via1 >>
rect 5690 12724 5742 12776
rect 5690 12660 5742 12712
rect 5819 12655 5871 12664
rect 5819 12621 5823 12655
rect 5823 12621 5857 12655
rect 5857 12621 5871 12655
rect 5819 12612 5871 12621
rect 5883 12655 5935 12664
rect 5883 12621 5895 12655
rect 5895 12621 5929 12655
rect 5929 12621 5935 12655
rect 5883 12612 5935 12621
rect 5690 12177 5742 12181
rect 5690 12143 5700 12177
rect 5700 12143 5734 12177
rect 5734 12143 5742 12177
rect 5690 12129 5742 12143
rect 5690 12105 5742 12117
rect 5690 12071 5700 12105
rect 5700 12071 5734 12105
rect 5734 12071 5742 12105
rect 5690 12065 5742 12071
rect 5688 10809 5740 10840
rect 5688 10788 5700 10809
rect 5700 10788 5734 10809
rect 5734 10788 5740 10809
rect 5688 10775 5700 10776
rect 5700 10775 5734 10776
rect 5734 10775 5740 10776
rect 5688 10729 5740 10775
rect 5688 10724 5700 10729
rect 5700 10724 5734 10729
rect 5734 10724 5740 10729
rect 5688 10615 5740 10622
rect 5688 10581 5700 10615
rect 5700 10581 5734 10615
rect 5734 10581 5740 10615
rect 5688 10570 5740 10581
rect 5688 10536 5740 10558
rect 5688 10506 5700 10536
rect 5700 10506 5734 10536
rect 5734 10506 5740 10536
rect 6154 12668 6206 12720
rect 6154 12604 6206 12656
rect 6069 10788 6121 10840
rect 6069 10724 6121 10776
rect 5847 9980 5899 10032
rect 5911 9980 5963 10032
rect 5975 9980 6027 10032
rect 5847 9898 5899 9950
rect 5911 9898 5963 9950
rect 5975 9898 6027 9950
rect 5847 9816 5899 9868
rect 5911 9816 5963 9868
rect 5975 9816 6027 9868
rect 5847 9733 5899 9785
rect 5911 9733 5963 9785
rect 5975 9733 6027 9785
rect 6154 10570 6206 10622
rect 6154 10506 6206 10558
rect 6069 9563 6121 9615
rect 6069 9499 6121 9551
rect 5704 9376 5756 9428
rect 5704 9312 5756 9364
rect 6066 9423 6118 9428
rect 6066 9389 6075 9423
rect 6075 9389 6109 9423
rect 6109 9389 6118 9423
rect 6066 9376 6118 9389
rect 6066 9312 6118 9364
rect 6157 9387 6209 9439
rect 6157 9323 6209 9375
rect -10457 8061 -10405 8113
rect -10391 8061 -10339 8113
rect -9494 8055 -9442 8107
rect 5430 8101 5482 8153
rect 5494 8101 5546 8153
rect 5931 9030 5983 9082
rect -9696 7996 -9644 8002
rect -9696 7962 -9687 7996
rect -9687 7962 -9653 7996
rect -9653 7962 -9644 7996
rect -9494 7989 -9442 8041
rect 5514 8017 5566 8069
rect 5578 8017 5630 8069
rect 5684 8953 5736 9005
rect 5684 8889 5736 8941
rect -9696 7950 -9644 7962
rect -9696 7924 -9644 7936
rect -9696 7890 -9687 7924
rect -9687 7890 -9653 7924
rect -9653 7890 -9644 7924
rect -9696 7884 -9644 7890
rect -9999 7807 -9947 7859
rect -9999 7741 -9947 7793
rect -9919 7712 -9910 7738
rect -9910 7712 -9876 7738
rect -9876 7712 -9867 7738
rect -9919 7686 -9867 7712
rect -9919 7663 -9867 7672
rect -10095 7589 -10043 7631
rect -9919 7629 -9910 7663
rect -9910 7629 -9876 7663
rect -9876 7629 -9867 7663
rect -9919 7620 -9867 7629
rect -9574 7734 -9568 7738
rect -9568 7734 -9534 7738
rect -9534 7734 -9522 7738
rect -9574 7687 -9522 7734
rect -9574 7686 -9568 7687
rect -9568 7686 -9534 7687
rect -9534 7686 -9522 7687
rect -9574 7653 -9568 7672
rect -9568 7653 -9534 7672
rect -9534 7653 -9522 7672
rect -9574 7620 -9522 7653
rect -10095 7579 -10086 7589
rect -10086 7579 -10052 7589
rect -10052 7579 -10043 7589
rect -10095 7555 -10086 7567
rect -10086 7555 -10052 7567
rect -10052 7555 -10043 7567
rect -10095 7515 -10043 7555
rect -10505 7455 -10453 7461
rect -10505 7421 -10490 7455
rect -10490 7421 -10456 7455
rect -10456 7421 -10453 7455
rect -10505 7409 -10453 7421
rect -9696 7572 -9644 7578
rect -9696 7538 -9687 7572
rect -9687 7538 -9653 7572
rect -9653 7538 -9644 7572
rect -9696 7526 -9644 7538
rect -9696 7500 -9644 7512
rect -9696 7466 -9687 7500
rect -9687 7466 -9653 7500
rect -9653 7466 -9644 7500
rect -9696 7460 -9644 7466
rect -9574 7444 -9522 7451
rect -9574 7410 -9568 7444
rect -9568 7410 -9534 7444
rect -9534 7410 -9522 7444
rect -9574 7399 -9522 7410
rect -10505 7383 -10453 7397
rect -10505 7349 -10490 7383
rect -10490 7349 -10456 7383
rect -10456 7349 -10453 7383
rect -10505 7345 -10453 7349
rect -10225 7353 -10173 7359
rect -10225 7319 -10219 7353
rect -10219 7319 -10185 7353
rect -10185 7319 -10173 7353
rect -10225 7307 -10173 7319
rect -10161 7353 -10109 7359
rect -10161 7319 -10147 7353
rect -10147 7319 -10113 7353
rect -10113 7319 -10109 7353
rect -10161 7307 -10109 7319
rect -10035 7365 -9983 7371
rect -10035 7331 -10029 7365
rect -10029 7331 -9995 7365
rect -9995 7331 -9983 7365
rect -10035 7319 -9983 7331
rect -9969 7365 -9917 7371
rect -9969 7331 -9957 7365
rect -9957 7331 -9923 7365
rect -9923 7331 -9917 7365
rect -9969 7319 -9917 7331
rect -9574 7363 -9522 7385
rect -9686 7280 -9634 7332
rect -9574 7333 -9568 7363
rect -9568 7333 -9534 7363
rect -9534 7333 -9522 7363
rect -9686 7214 -9634 7266
rect 5598 7933 5650 7985
rect 5662 7933 5714 7985
rect 5681 7849 5733 7901
rect 5745 7849 5797 7901
rect 5848 8927 5900 8979
rect 5848 8863 5900 8915
rect 5761 7765 5813 7817
rect 5825 7765 5877 7817
rect 5931 8966 5983 9018
rect 5861 7681 5913 7733
rect 5925 7681 5977 7733
rect 6025 8895 6077 8947
rect 6025 8831 6077 8883
rect 5955 7597 6007 7649
rect 6019 7597 6071 7649
rect 6066 7513 6118 7565
rect 6130 7513 6182 7565
rect -9494 7113 -9442 7165
rect -9494 7047 -9442 7099
rect -10459 6714 -10447 6748
rect -10447 6714 -10413 6748
rect -10413 6714 -10407 6748
rect -10459 6696 -10407 6714
rect -10459 6627 -10407 6679
rect -10459 6558 -10407 6610
rect -9971 6416 -9919 6468
rect -9898 6416 -9846 6468
rect -9233 6406 -9181 6458
rect -9160 6406 -9108 6458
rect -9971 6370 -9919 6382
rect -9971 6336 -9967 6370
rect -9967 6336 -9933 6370
rect -9933 6336 -9919 6370
rect -9971 6330 -9919 6336
rect -9898 6370 -9846 6382
rect -9898 6336 -9886 6370
rect -9886 6336 -9852 6370
rect -9852 6336 -9846 6370
rect -9898 6330 -9846 6336
rect -9664 6370 -9612 6376
rect -9591 6370 -9539 6376
rect -9664 6336 -9657 6370
rect -9657 6336 -9618 6370
rect -9618 6336 -9612 6370
rect -9591 6336 -9584 6370
rect -9584 6336 -9545 6370
rect -9545 6336 -9539 6370
rect -9664 6324 -9612 6336
rect -9591 6324 -9539 6336
rect -8041 6370 -7989 6376
rect -8041 6336 -8035 6370
rect -8035 6336 -8001 6370
rect -8001 6336 -7989 6370
rect -8041 6324 -7989 6336
rect -7968 6370 -7916 6376
rect -7968 6336 -7961 6370
rect -7961 6336 -7927 6370
rect -7927 6336 -7916 6370
rect -7968 6324 -7916 6336
rect -6186 6370 -6134 6376
rect -6113 6370 -6061 6376
rect -6186 6336 -6160 6370
rect -6160 6336 -6134 6370
rect -6113 6336 -6087 6370
rect -6087 6336 -6061 6370
rect -6186 6324 -6134 6336
rect -6113 6324 -6061 6336
rect -5553 6296 -5501 6348
rect -5489 6296 -5437 6348
rect -3730 6235 -3678 6287
rect -3666 6235 -3614 6287
rect -9233 6171 -9181 6223
rect -9160 6171 -9108 6223
rect -8041 6171 -7989 6223
rect -7968 6171 -7916 6223
rect -10459 6104 -10407 6156
rect -10459 6035 -10407 6087
rect -10459 5966 -10407 6018
rect -9977 6079 -9925 6131
rect -9800 6110 -9748 6162
rect -9727 6110 -9675 6162
rect -9977 6014 -9925 6066
rect -6886 6008 -6834 6060
rect -6817 6008 -6765 6060
rect -6748 6008 -6696 6060
rect -5365 6051 -5313 6103
rect -5292 6051 -5240 6103
rect -5219 6051 -5167 6103
rect -5146 6051 -5094 6103
<< metal2 >>
rect 5690 12776 5742 12782
rect 5690 12712 5742 12724
rect 6154 12720 6206 12726
rect 6154 12664 6206 12668
rect 5690 12181 5742 12660
rect 5813 12612 5819 12664
rect 5871 12612 5883 12664
rect 5935 12656 6206 12664
rect 5935 12612 6154 12656
rect 5938 12611 6154 12612
rect 6154 12598 6206 12604
rect 5690 12117 5742 12129
rect 5690 12059 5742 12065
rect 5688 10840 6121 10846
rect 5740 10788 6069 10840
rect 5688 10776 6121 10788
rect 5740 10724 6069 10776
rect 5688 10718 6121 10724
rect 5688 10622 6206 10628
rect 5740 10570 6154 10622
rect 5688 10558 6206 10570
rect 5740 10506 6154 10558
rect 5688 10500 6206 10506
rect 5846 10032 6028 10038
rect 5846 9972 5847 10032
rect 5899 10028 5911 10032
rect 5903 9980 5911 10028
rect 5963 10028 5975 10032
rect 5963 9980 5971 10028
rect 5903 9972 5971 9980
rect 6027 9972 6028 10032
rect 5846 9950 6028 9972
rect 5846 9816 5847 9950
rect 5899 9911 5911 9950
rect 5903 9898 5911 9911
rect 5963 9911 5975 9950
rect 5963 9898 5971 9911
rect 5903 9868 5971 9898
rect 5903 9855 5911 9868
rect 5899 9816 5911 9855
rect 5963 9855 5971 9868
rect 5963 9816 5975 9855
rect 6027 9816 6028 9950
rect 5846 9793 6028 9816
rect 5846 9733 5847 9793
rect 5903 9785 5971 9793
rect 5903 9737 5911 9785
rect 5899 9733 5911 9737
rect 5963 9737 5971 9785
rect 5963 9733 5975 9737
rect 6027 9733 6028 9793
rect 5846 9727 6028 9733
rect 5617 9615 6121 9621
rect 5617 9563 6069 9615
rect 5617 9551 6121 9563
rect 5617 9499 6069 9551
rect 5617 9493 6121 9499
rect 5617 9032 5669 9493
rect 6157 9439 6209 9445
rect 5704 9428 5756 9434
tri 5756 9428 5762 9434 sw
rect 6066 9428 6118 9434
rect 5756 9389 5762 9428
tri 5762 9389 5801 9428 sw
rect 5756 9376 6066 9389
rect 5704 9364 6118 9376
rect 5756 9312 6066 9364
rect 5704 9306 6118 9312
rect 6157 9375 6209 9387
tri 6122 9088 6157 9123 se
rect 6157 9088 6209 9323
rect 5931 9082 6209 9088
tri 5669 9032 5715 9078 sw
rect 5617 9030 5715 9032
tri 5715 9030 5717 9032 sw
rect 5983 9030 6209 9082
rect 5617 9029 5717 9030
tri 5717 9029 5718 9030 sw
tri 5617 9018 5628 9029 ne
rect 5628 9018 5718 9029
tri 5718 9018 5729 9029 sw
rect 5931 9026 6209 9030
rect 5931 9018 5983 9026
tri 5628 9011 5635 9018 ne
rect 5635 9011 5729 9018
tri 5729 9011 5736 9018 sw
tri 5635 9005 5641 9011 ne
rect 5641 9005 5736 9011
tri 5641 8962 5684 9005 ne
rect 5684 8941 5736 8953
rect 5684 8883 5736 8889
rect 5848 8979 5900 8985
tri 5983 8990 6019 9026 nw
rect 5931 8960 5983 8966
rect 5848 8915 5900 8927
rect 6025 8947 6077 8953
rect 5848 8857 5900 8863
rect 5957 8860 5966 8916
rect 6022 8895 6025 8916
rect 6022 8883 6046 8895
rect 6022 8860 6025 8883
rect 6102 8860 6111 8916
tri 5991 8857 5994 8860 ne
rect 5994 8857 6025 8860
tri 5994 8831 6020 8857 ne
rect 6020 8831 6025 8857
tri 6020 8826 6025 8831 ne
rect 6025 8825 6077 8831
tri 6077 8826 6111 8860 nw
tri 4738 8140 4751 8153 se
rect 4751 8140 5430 8153
rect -10463 8061 -10457 8113
rect -10405 8061 -10391 8113
rect -10339 8107 -9442 8113
rect -10339 8061 -9494 8107
tri -9530 8055 -9524 8061 ne
rect -9524 8055 -9494 8061
tri -9524 8041 -9510 8055 ne
rect -9510 8041 -9442 8055
tri -9510 8025 -9494 8041 ne
tri -10043 8003 -10038 8008 se
rect -10038 8003 -9644 8008
tri -10044 8002 -10043 8003 se
rect -10043 8002 -9644 8003
tri -10094 7952 -10044 8002 se
rect -10044 7952 -9696 8002
tri -10095 7951 -10094 7952 se
rect -10094 7951 -10014 7952
rect -10095 7950 -10014 7951
tri -10014 7950 -10012 7952 nw
tri -9731 7950 -9729 7952 ne
rect -9729 7950 -9696 7952
rect -9494 7983 -9442 7989
rect 4738 8101 5430 8140
rect 5482 8101 5494 8153
rect 5546 8101 5569 8153
rect -10095 7936 -10028 7950
tri -10028 7936 -10014 7950 nw
tri -9729 7936 -9715 7950 ne
rect -9715 7936 -9644 7950
rect -10095 7631 -10043 7936
tri -10043 7921 -10028 7936 nw
tri -9715 7921 -9700 7936 ne
rect -9700 7921 -9696 7936
tri -9700 7917 -9696 7921 ne
rect -9696 7878 -9644 7884
rect -10095 7567 -10043 7579
rect -10095 7509 -10043 7515
rect -9999 7859 -9947 7865
rect -9999 7793 -9947 7807
rect -9999 7597 -9947 7741
rect -9919 7738 -9867 7744
rect -9574 7738 -9522 7744
tri -9867 7692 -9841 7718 sw
tri -9600 7692 -9574 7718 se
rect -9867 7686 -9574 7692
rect -9919 7672 -9522 7686
rect -9867 7640 -9574 7672
rect -9867 7620 -9861 7640
tri -9861 7620 -9841 7640 nw
tri -9600 7620 -9580 7640 ne
rect -9580 7620 -9574 7640
rect -9919 7614 -9867 7620
tri -9867 7614 -9861 7620 nw
tri -9580 7614 -9574 7620 ne
rect -9574 7614 -9522 7620
tri -9947 7597 -9942 7602 sw
rect -9999 7578 -9942 7597
tri -9942 7578 -9923 7597 sw
rect -9696 7578 -9644 7584
rect -9999 7567 -9923 7578
tri -9923 7567 -9912 7578 sw
rect -9999 7507 -9754 7567
tri -9857 7488 -9838 7507 ne
rect -9838 7488 -9754 7507
tri -9838 7467 -9817 7488 ne
rect -9817 7467 -9754 7488
rect -10505 7461 -10453 7467
tri -9817 7460 -9810 7467 ne
rect -9810 7460 -9754 7467
tri -9810 7456 -9806 7460 ne
rect -10505 7397 -10453 7409
rect -10505 6756 -10453 7345
rect -10231 7307 -10225 7359
rect -10173 7307 -10161 7359
rect -10109 7307 -10103 7359
rect -10041 7319 -10035 7371
rect -9983 7319 -9969 7371
rect -9917 7319 -9911 7371
tri -10019 7307 -10007 7319 ne
rect -10007 7307 -9925 7319
tri -9925 7307 -9913 7319 nw
tri -10007 7280 -9980 7307 ne
rect -9980 7280 -9925 7307
tri -9980 7277 -9977 7280 ne
tri -10505 6754 -10503 6756 ne
rect -10503 6754 -10453 6756
tri -10453 6754 -10407 6800 sw
tri -10503 6748 -10497 6754 ne
rect -10497 6748 -10407 6754
tri -10497 6710 -10459 6748 ne
rect -10459 6679 -10407 6696
rect -10459 6610 -10407 6627
rect -10459 6156 -10407 6558
rect -9977 6468 -9925 7280
rect -9977 6416 -9971 6468
rect -9919 6416 -9898 6468
rect -9846 6416 -9840 6468
rect -10459 6087 -10407 6104
rect -10459 6018 -10407 6035
rect -9977 6330 -9971 6382
rect -9919 6330 -9898 6382
rect -9846 6330 -9840 6382
rect -9977 6131 -9925 6330
rect -9806 6171 -9754 7460
rect -9644 7526 -9162 7540
rect -9696 7512 -9162 7526
rect -9644 7488 -9162 7512
rect -9696 7454 -9644 7460
rect -9574 7451 -9522 7457
tri -9522 7405 -9496 7431 sw
rect -9522 7399 -9262 7405
rect -9574 7385 -9262 7399
rect -9686 7332 -9634 7338
rect -9522 7353 -9262 7385
rect -9522 7338 -9511 7353
tri -9511 7338 -9496 7353 nw
rect -9574 7327 -9522 7333
tri -9522 7327 -9511 7338 nw
rect -9686 7266 -9634 7280
rect -9686 6955 -9634 7214
rect -9314 7177 -9262 7353
rect -9214 7265 -9162 7488
rect -9214 7213 -7714 7265
rect -9494 7165 -9442 7171
rect -9314 7154 -7819 7177
tri -7819 7154 -7796 7177 sw
rect -9314 7125 -7796 7154
rect -9494 7099 -9442 7113
tri -7878 7095 -7848 7125 ne
rect -9442 7064 -7907 7093
tri -7907 7064 -7878 7093 sw
rect -9442 7047 -7878 7064
rect -9494 7041 -7878 7047
tri -9686 6907 -9638 6955 ne
rect -9638 6907 -9634 6955
tri -9634 6907 -9559 6982 sw
tri -9638 6903 -9634 6907 ne
rect -9634 6903 -9559 6907
tri -9634 6876 -9607 6903 ne
tri -9612 6406 -9607 6411 se
rect -9607 6406 -9559 6903
rect -7921 6458 -7878 7041
rect -7848 6539 -7796 7125
rect -7766 6619 -7714 7213
tri -7714 6619 -7680 6653 sw
rect -7766 6601 -2300 6619
tri -7766 6567 -7732 6601 ne
rect -7732 6567 -2300 6601
rect -7848 6487 -2397 6539
tri -7878 6458 -7863 6473 sw
tri -9614 6404 -9612 6406 se
rect -9612 6404 -9559 6406
tri -9616 6402 -9614 6404 se
rect -9614 6402 -9559 6404
rect -9239 6406 -9233 6458
rect -9181 6406 -9160 6458
rect -9108 6406 -9102 6458
rect -7921 6450 -7863 6458
tri -7863 6450 -7855 6458 sw
rect -7921 6424 -3803 6450
tri -3803 6424 -3777 6450 sw
rect -7921 6423 -3777 6424
tri -7921 6406 -7904 6423 ne
rect -7904 6406 -3777 6423
tri -9636 6382 -9616 6402 se
rect -9616 6382 -9559 6402
tri -9559 6382 -9539 6402 sw
tri -9642 6376 -9636 6382 se
rect -9636 6376 -9539 6382
tri -9539 6376 -9533 6382 sw
rect -9670 6324 -9664 6376
rect -9612 6324 -9591 6376
rect -9539 6324 -9533 6376
rect -9239 6223 -9102 6406
tri -7904 6404 -7902 6406 ne
rect -7902 6404 -3777 6406
tri -3871 6382 -3849 6404 ne
rect -3849 6382 -3777 6404
tri -3849 6376 -3843 6382 ne
rect -3843 6376 -3777 6382
tri -9754 6171 -9731 6194 sw
rect -9239 6171 -9233 6223
rect -9181 6171 -9160 6223
rect -9108 6171 -9102 6223
rect -8047 6324 -8041 6376
rect -7989 6324 -7968 6376
rect -7916 6324 -7910 6376
rect -8047 6223 -7910 6324
rect -8047 6171 -8041 6223
rect -7989 6171 -7968 6223
rect -7916 6171 -7910 6223
rect -6192 6324 -6186 6376
rect -6134 6324 -6113 6376
rect -6061 6324 -6055 6376
tri -3843 6359 -3826 6376 ne
rect -9806 6162 -9731 6171
tri -9731 6162 -9722 6171 sw
rect -9806 6110 -9800 6162
rect -9748 6110 -9727 6162
rect -9675 6110 -9669 6162
rect -9977 6066 -9925 6079
rect -9977 6008 -9925 6014
rect -6892 6008 -6886 6060
rect -6834 6008 -6817 6060
rect -6765 6008 -6748 6060
rect -6696 6051 -6582 6060
tri -6582 6051 -6573 6060 sw
rect -6696 6008 -6573 6051
tri -6573 6008 -6530 6051 sw
rect -10459 5960 -10407 5966
tri -6612 5960 -6564 6008 ne
rect -6564 5960 -6530 6008
tri -6564 5939 -6543 5960 ne
rect -6543 5939 -6530 5960
tri -6530 5939 -6461 6008 sw
tri -6543 5867 -6471 5939 ne
rect -6471 5867 -6461 5939
tri -6461 5867 -6389 5939 sw
rect -6192 5919 -6055 6324
rect -5559 6296 -5553 6348
rect -5501 6296 -5489 6348
rect -5437 6296 -5431 6348
rect -5559 6011 -5431 6296
rect -3826 6195 -3777 6376
rect -2449 6383 -2397 6487
rect -2352 6463 -2300 6567
tri 4703 6466 4738 6501 se
rect 4738 6467 4790 8101
rect 4738 6466 4789 6467
tri 4789 6466 4790 6467 nw
tri 4822 8056 4835 8069 se
rect 4835 8056 5514 8069
rect 4822 8017 5514 8056
rect 5566 8017 5578 8069
rect 5630 8017 5636 8069
tri 4700 6463 4703 6466 se
rect 4703 6463 4786 6466
tri 4786 6463 4789 6466 nw
rect -2352 6429 4752 6463
tri 4752 6429 4786 6463 nw
rect -2352 6411 4734 6429
tri 4734 6411 4752 6429 nw
tri 4804 6411 4822 6429 se
rect 4822 6411 4874 8017
tri 4776 6383 4804 6411 se
rect 4804 6402 4874 6411
rect 4804 6383 4855 6402
tri 4855 6383 4874 6402 nw
tri 4906 7961 4930 7985 se
rect 4930 7961 5598 7985
rect 4906 7933 5598 7961
rect 5650 7933 5662 7985
rect 5714 7933 5720 7985
rect -2449 6331 4803 6383
tri 4803 6331 4855 6383 nw
rect 4906 6287 4958 7933
rect -3736 6235 -3730 6287
rect -3678 6235 -3666 6287
rect -3614 6235 4958 6287
tri 4990 7882 5009 7901 se
rect 5009 7882 5681 7901
rect 4990 7849 5681 7882
rect 5733 7849 5745 7901
rect 5797 7849 5803 7901
tri -3777 6195 -3746 6226 sw
rect 4990 6195 5042 7849
rect -3826 6143 5042 6195
tri 5074 7803 5088 7817 se
rect 5088 7803 5761 7817
rect 5074 7765 5761 7803
rect 5813 7765 5825 7817
rect 5877 7765 5883 7817
rect 5074 6103 5126 7765
rect -5371 6051 -5365 6103
rect -5313 6051 -5292 6103
rect -5240 6051 -5219 6103
rect -5167 6051 -5146 6103
rect -5094 6051 5126 6103
tri 5158 7709 5182 7733 se
rect 5182 7709 5861 7733
rect 5158 7681 5861 7709
rect 5913 7681 5925 7733
rect 5977 7681 5983 7733
rect 5158 6011 5210 7681
rect -5559 5959 5210 6011
tri 5242 7630 5261 7649 se
rect 5261 7630 5955 7649
rect 5242 7597 5955 7630
rect 6007 7597 6019 7649
rect 6071 7597 6077 7649
rect 5242 5919 5294 7597
rect -6192 5867 5294 5919
tri 5326 7545 5346 7565 se
rect 5346 7545 6066 7565
rect 5326 7513 6066 7545
rect 6118 7513 6130 7565
rect 6182 7513 6188 7565
tri -6471 5857 -6461 5867 ne
rect -6461 5857 -6389 5867
tri -6389 5857 -6379 5867 sw
tri -6461 5827 -6431 5857 ne
rect -6431 5827 -6379 5857
tri -6379 5827 -6349 5857 sw
rect 5326 5827 5378 7513
tri -6431 5775 -6379 5827 ne
rect -6379 5775 5378 5827
<< via2 >>
rect 5847 9980 5899 10028
rect 5899 9980 5903 10028
rect 5971 9980 5975 10028
rect 5975 9980 6027 10028
rect 5847 9972 5903 9980
rect 5971 9972 6027 9980
rect 5847 9898 5899 9911
rect 5899 9898 5903 9911
rect 5971 9898 5975 9911
rect 5975 9898 6027 9911
rect 5847 9868 5903 9898
rect 5971 9868 6027 9898
rect 5847 9855 5899 9868
rect 5899 9855 5903 9868
rect 5971 9855 5975 9868
rect 5975 9855 6027 9868
rect 5847 9785 5903 9793
rect 5971 9785 6027 9793
rect 5847 9737 5899 9785
rect 5899 9737 5903 9785
rect 5971 9737 5975 9785
rect 5975 9737 6027 9785
rect 5966 8860 6022 8916
rect 6046 8895 6077 8916
rect 6077 8895 6102 8916
rect 6046 8883 6102 8895
rect 6046 8860 6077 8883
rect 6077 8860 6102 8883
<< metal3 >>
rect 5842 10028 6032 10033
rect 5842 9972 5847 10028
rect 5903 9972 5971 10028
rect 6027 9972 6032 10028
rect 5842 9911 6032 9972
rect 5842 9855 5847 9911
rect 5903 9855 5971 9911
rect 6027 9855 6032 9911
rect 5842 9793 6032 9855
rect 5842 9737 5847 9793
rect 5903 9737 5971 9793
rect 6027 9737 6032 9793
rect 5842 9732 6032 9737
rect 5961 8916 6107 8921
rect 5961 8860 5966 8916
rect 6022 8860 6046 8916
rect 6102 8860 6107 8916
rect 5961 8855 6107 8860
use sky130_fd_pr__nfet_01v8__example_5595914180817  sky130_fd_pr__nfet_01v8__example_5595914180817_0
timestamp 1663361622
transform 1 0 -10294 0 1 5964
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180818  sky130_fd_pr__nfet_01v8__example_5595914180818_0
timestamp 1663361622
transform -1 0 -9921 0 -1 8001
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180818  sky130_fd_pr__nfet_01v8__example_5595914180818_1
timestamp 1663361622
transform -1 0 -10097 0 -1 8001
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180865  sky130_fd_pr__nfet_01v8__example_5595914180865_0
timestamp 1663361622
transform -1 0 -6447 0 -1 6618
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_5595914180865  sky130_fd_pr__nfet_01v8__example_5595914180865_1
timestamp 1663361622
transform -1 0 -8103 0 -1 6618
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_5595914180866  sky130_fd_pr__nfet_01v8__example_5595914180866_0
timestamp 1663361622
transform -1 0 -9759 0 -1 6618
box -1 0 801 1
use sky130_fd_pr__nfet_01v8__example_5595914180866  sky130_fd_pr__nfet_01v8__example_5595914180866_1
timestamp 1663361622
transform -1 0 -5591 0 -1 6618
box -1 0 801 1
use sky130_fd_pr__nfet_01v8__example_5595914180867  sky130_fd_pr__nfet_01v8__example_5595914180867_0
timestamp 1663361622
transform 0 -1 -9616 1 0 7086
box -1 0 857 1
use sky130_fd_pr__nfet_01v8__example_5595914180870  sky130_fd_pr__nfet_01v8__example_5595914180870_0
timestamp 1663361622
transform 0 -1 -10432 1 0 7457
box -1 0 401 1
use sky130_fd_pr__pfet_01v8__example_5595914180871  sky130_fd_pr__pfet_01v8__example_5595914180871_0
timestamp 1663361622
transform 1 0 5821 0 1 12433
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_5595914180871  sky130_fd_pr__pfet_01v8__example_5595914180871_1
timestamp 1663361622
transform 1 0 6179 0 1 12433
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_5595914180873  sky130_fd_pr__pfet_01v8__example_5595914180873_0
timestamp 1663361622
transform 0 -1 6382 1 0 12059
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_5595914180874  sky130_fd_pr__pfet_01v8__example_5595914180874_0
timestamp 1663361622
transform 1 0 5958 0 -1 9432
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_5595914180876  sky130_fd_pr__pfet_01v8__example_5595914180876_0
timestamp 1663361622
transform 0 -1 6382 1 0 10683
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_5595914180876  sky130_fd_pr__pfet_01v8__example_5595914180876_1
timestamp 1663361622
transform 0 -1 6382 1 0 9659
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_5595914180876  sky130_fd_pr__pfet_01v8__example_5595914180876_2
timestamp 1663361622
transform 0 -1 6382 1 0 10171
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_5595914180876  sky130_fd_pr__pfet_01v8__example_5595914180876_3
timestamp 1663361622
transform 0 -1 6382 1 0 11195
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_5595914180877  sky130_fd_pr__pfet_01v8__example_5595914180877_0
timestamp 1663361622
transform 0 -1 6382 1 0 11707
box -1 0 297 1
<< labels >>
flabel metal1 s 5918 11773 6031 11926 0 FreeSans 600 0 0 0 VPWR
port 1 nsew
flabel metal1 s -10458 6559 -10288 6657 3 FreeSans 520 180 0 0 VGND
port 2 nsew
flabel metal1 s -10373 6608 -10373 6608 3 FreeSans 520 180 0 0 VGND
port 2 nsew
flabel comment s 6293 11866 6293 11866 0 FreeSans 200 270 0 0 P1G
flabel comment s 5778 11848 5778 11848 0 FreeSans 200 90 0 0 P1GB
flabel comment s 5937 12634 5937 12634 0 FreeSans 200 180 0 0 P1G_NEW
flabel comment s 6215 12492 6215 12492 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6034 12492 6034 12492 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6389 12504 6389 12504 0 FreeSans 200 90 0 0 P2GB
flabel comment s 5852 12504 5852 12504 0 FreeSans 200 90 0 0 P1GB
flabel comment s 6119 10657 6119 10657 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6119 10142 6119 10142 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6119 9633 6119 9633 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6160 10404 6160 10404 0 FreeSans 200 90 0 0 P2G_NEW
flabel comment s 6160 9887 6160 9887 0 FreeSans 200 90 0 0 P2G_NEW
flabel comment s 5779 11428 5779 11428 0 FreeSans 200 90 0 0 PADLO
flabel comment s 5778 10911 5778 10911 0 FreeSans 200 90 0 0 P2G_NEW
flabel comment s 5778 9887 5778 9887 0 FreeSans 200 90 0 0 PADLO_BAR
flabel comment s 5779 10404 5779 10404 0 FreeSans 200 90 0 0 P1G_NEW
flabel comment s 6160 9168 6160 9168 0 FreeSans 200 180 0 0 PADLO
flabel comment s 5778 12125 5778 12125 0 FreeSans 200 90 0 0 P2GB
flabel comment s 6089 12031 6089 12031 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6089 11675 6089 11675 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6293 12207 6293 12207 0 FreeSans 200 270 0 0 P2G
flabel comment s 6169 9333 6169 9333 0 FreeSans 200 90 0 0 PADLO_BAR
flabel comment s 5991 9316 5991 9316 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6343 9316 6343 9316 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6298 12634 6298 12634 0 FreeSans 200 180 0 0 P2G_NEW
flabel comment s 6119 10657 6119 10657 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6119 11166 6119 11166 0 FreeSans 200 90 0 0 VPWR
flabel comment s 6241 11428 6241 11428 0 FreeSans 200 90 0 0 P1G_NEW
flabel comment s 6247 10911 6247 10911 0 FreeSans 200 90 0 0 P1G_NEW
flabel comment s -1754 5913 -1754 5913 0 FreeSans 400 0 0 0 PADLO
flabel comment s -1754 6002 -1754 6002 0 FreeSans 400 0 0 0 P1G_NEW
flabel comment s -1754 6271 -1754 6271 0 FreeSans 400 0 0 0 P2G_NEW
flabel comment s -1754 6090 -1754 6090 0 FreeSans 400 0 0 0 P1GB
flabel comment s -8071 6556 -8071 6556 0 FreeSans 400 270 0 0 VGND
flabel comment s -10081 6663 -10081 6663 0 FreeSans 400 270 0 0 VGND
flabel comment s -1754 6182 -1754 6182 0 FreeSans 400 0 0 0 P1G
flabel comment s -1754 6371 -1754 6371 0 FreeSans 400 0 0 0 P2GB
flabel comment s -169 5972 -169 5972 0 FreeSans 200 0 0 0 P2G
flabel comment s 5855 9215 5855 9215 0 FreeSans 200 270 0 0 PADLO
flabel comment s 5777 9271 5777 9271 0 FreeSans 200 90 0 0 PADLO_BAR
flabel comment s 5557 9069 5557 9069 0 FreeSans 200 270 0 0 P2G
flabel comment s 6338 9069 6338 9069 0 FreeSans 200 270 0 0 P1G
flabel comment s 6247 9112 6247 9112 0 FreeSans 200 90 0 0 P1G_NEW
flabel comment s 6408 9080 6408 9080 0 FreeSans 200 90 0 0 P2GB
flabel comment s 5698 9024 5698 9024 0 FreeSans 200 90 0 0 P2G_NEW
flabel comment s -1754 6450 -1754 6450 0 FreeSans 400 0 0 0 P2G
flabel comment s -1754 5816 -1754 5816 0 FreeSans 400 0 0 0 PADLO_BAR
flabel comment s 5391 8126 5391 8126 0 FreeSans 200 0 0 0 P2G
flabel comment s 5683 9199 5683 9199 0 FreeSans 200 90 0 0 P1GB
flabel comment s -922 5913 -922 5913 0 FreeSans 400 0 0 0 PADLO
flabel comment s -922 6002 -922 6002 0 FreeSans 400 0 0 0 P1G_NEW
flabel comment s -922 6090 -922 6090 0 FreeSans 400 0 0 0 P1GB
flabel comment s -922 6371 -922 6371 0 FreeSans 400 0 0 0 P2GB
flabel comment s -922 6182 -922 6182 0 FreeSans 400 0 0 0 P1G
flabel comment s -922 6450 -922 6450 0 FreeSans 400 0 0 0 P2G
flabel comment s -922 6271 -922 6271 0 FreeSans 400 0 0 0 P2G_NEW
flabel comment s -922 5816 -922 5816 0 FreeSans 400 0 0 0 PADLO_BAR
flabel comment s 6144 8126 6144 8126 0 FreeSans 400 270 0 0 PADLO_BAR
flabel comment s 4929 6768 4929 6768 0 FreeSans 400 90 0 0 P2G_NEW
flabel comment s 4759 6768 4759 6768 0 FreeSans 400 90 0 0 P2G
flabel comment s 5018 6768 5018 6768 0 FreeSans 400 90 0 0 P1G
flabel comment s 4838 6768 4838 6768 0 FreeSans 400 90 0 0 P2GB
flabel comment s 5094 6768 5094 6768 0 FreeSans 400 90 0 0 P1GB
flabel comment s 5182 6768 5182 6768 0 FreeSans 400 90 0 0 P1G_NEW
flabel comment s 5271 6768 5271 6768 0 FreeSans 400 90 0 0 PADLO
flabel comment s 5348 6757 5348 6757 0 FreeSans 400 90 0 0 PADLO_BAR
flabel metal2 s 4990 7506 5042 7565 0 FreeSans 200 0 0 0 P1G
port 3 nsew
flabel metal2 s 5244 7510 5293 7562 0 FreeSans 200 0 0 0 PADLO
port 4 nsew
flabel metal2 s 5723 7779 5750 7806 0 FreeSans 200 0 0 0 P1GB
port 5 nsew
flabel metal2 s -1651 6411 -1599 6463 0 FreeSans 200 0 0 0 P2G
port 6 nsew
<< properties >>
string GDS_END 35412546
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 35321928
<< end >>
