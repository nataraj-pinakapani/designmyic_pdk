magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 4305 -208 4839 64
<< pwell >>
rect 72 1803 424 2217
rect 1105 2123 1357 2661
rect 1105 955 1590 2123
rect 1106 10 1590 955
rect 1504 2 1590 10
<< mvnmos >>
rect 98 2038 398 2138
rect 98 1882 398 1982
rect 1132 682 1432 782
rect 1132 526 1432 626
rect 1132 245 1432 345
rect 1132 89 1432 189
<< mvpmos >>
rect 4424 -142 4544 -2
rect 4600 -142 4720 -2
<< mvnnmos >>
rect 1131 1863 1331 2043
rect 1131 1627 1331 1807
rect 1131 1270 1331 1450
rect 1131 1034 1331 1214
<< nmoslvt >>
rect 1131 2552 1331 2582
rect 1131 2466 1331 2496
rect 1131 2380 1331 2410
rect 1131 2294 1331 2324
<< ndiff >>
rect 1131 2627 1331 2635
rect 1131 2593 1149 2627
rect 1183 2593 1217 2627
rect 1251 2593 1285 2627
rect 1319 2593 1331 2627
rect 1131 2582 1331 2593
rect 1131 2541 1331 2552
rect 1131 2507 1149 2541
rect 1183 2507 1217 2541
rect 1251 2507 1285 2541
rect 1319 2507 1331 2541
rect 1131 2496 1331 2507
rect 1131 2455 1331 2466
rect 1131 2421 1149 2455
rect 1183 2421 1217 2455
rect 1251 2421 1285 2455
rect 1319 2421 1331 2455
rect 1131 2410 1331 2421
rect 1131 2369 1331 2380
rect 1131 2335 1149 2369
rect 1183 2335 1217 2369
rect 1251 2335 1285 2369
rect 1319 2335 1331 2369
rect 1131 2324 1331 2335
rect 1131 2283 1331 2294
rect 1131 2249 1149 2283
rect 1183 2249 1217 2283
rect 1251 2249 1285 2283
rect 1319 2249 1331 2283
rect 1131 2241 1331 2249
<< mvndiff >>
rect 98 2183 398 2191
rect 98 2149 148 2183
rect 182 2149 216 2183
rect 250 2149 284 2183
rect 318 2149 352 2183
rect 386 2149 398 2183
rect 98 2138 398 2149
rect 1131 2088 1331 2096
rect 1131 2054 1149 2088
rect 1183 2054 1217 2088
rect 1251 2054 1285 2088
rect 1319 2054 1331 2088
rect 1131 2043 1331 2054
rect 98 2027 398 2038
rect 98 1993 148 2027
rect 182 1993 216 2027
rect 250 1993 284 2027
rect 318 1993 352 2027
rect 386 1993 398 2027
rect 98 1982 398 1993
rect 98 1871 398 1882
rect 98 1837 148 1871
rect 182 1837 216 1871
rect 250 1837 284 1871
rect 318 1837 352 1871
rect 386 1837 398 1871
rect 98 1829 398 1837
rect 1131 1852 1331 1863
rect 1131 1818 1149 1852
rect 1183 1818 1217 1852
rect 1251 1818 1285 1852
rect 1319 1818 1331 1852
rect 1131 1807 1331 1818
rect 1131 1616 1331 1627
rect 1131 1582 1149 1616
rect 1183 1582 1217 1616
rect 1251 1582 1285 1616
rect 1319 1582 1331 1616
rect 1131 1574 1331 1582
rect 1131 1495 1331 1503
rect 1131 1461 1143 1495
rect 1177 1461 1211 1495
rect 1245 1461 1279 1495
rect 1313 1461 1331 1495
rect 1131 1450 1331 1461
rect 1131 1259 1331 1270
rect 1131 1225 1143 1259
rect 1177 1225 1211 1259
rect 1245 1225 1279 1259
rect 1313 1225 1331 1259
rect 1131 1214 1331 1225
rect 1131 1023 1331 1034
rect 1131 989 1143 1023
rect 1177 989 1211 1023
rect 1245 989 1279 1023
rect 1313 989 1331 1023
rect 1131 981 1331 989
rect 1132 827 1432 835
rect 1132 793 1144 827
rect 1178 793 1212 827
rect 1246 793 1280 827
rect 1314 793 1348 827
rect 1382 793 1432 827
rect 1132 782 1432 793
rect 1132 671 1432 682
rect 1132 637 1144 671
rect 1178 637 1212 671
rect 1246 637 1280 671
rect 1314 637 1348 671
rect 1382 637 1432 671
rect 1132 626 1432 637
rect 1132 515 1432 526
rect 1132 481 1144 515
rect 1178 481 1212 515
rect 1246 481 1280 515
rect 1314 481 1348 515
rect 1382 481 1432 515
rect 1132 473 1432 481
rect 1132 390 1432 398
rect 1132 356 1144 390
rect 1178 356 1212 390
rect 1246 356 1280 390
rect 1314 356 1348 390
rect 1382 356 1432 390
rect 1132 345 1432 356
rect 1132 234 1432 245
rect 1132 200 1144 234
rect 1178 200 1212 234
rect 1246 200 1280 234
rect 1314 200 1348 234
rect 1382 200 1432 234
rect 1132 189 1432 200
rect 1132 78 1432 89
rect 1132 44 1144 78
rect 1178 44 1212 78
rect 1246 44 1280 78
rect 1314 44 1348 78
rect 1382 44 1432 78
rect 1132 36 1432 44
<< mvpdiff >>
rect 4371 -28 4424 -2
rect 4371 -62 4379 -28
rect 4413 -62 4424 -28
rect 4371 -96 4424 -62
rect 4371 -130 4379 -96
rect 4413 -130 4424 -96
rect 4371 -142 4424 -130
rect 4544 -28 4600 -2
rect 4544 -62 4555 -28
rect 4589 -62 4600 -28
rect 4544 -96 4600 -62
rect 4544 -130 4555 -96
rect 4589 -130 4600 -96
rect 4544 -142 4600 -130
rect 4720 -28 4773 -2
rect 4720 -62 4731 -28
rect 4765 -62 4773 -28
rect 4720 -96 4773 -62
rect 4720 -130 4731 -96
rect 4765 -130 4773 -96
rect 4720 -142 4773 -130
<< ndiffc >>
rect 1149 2593 1183 2627
rect 1217 2593 1251 2627
rect 1285 2593 1319 2627
rect 1149 2507 1183 2541
rect 1217 2507 1251 2541
rect 1285 2507 1319 2541
rect 1149 2421 1183 2455
rect 1217 2421 1251 2455
rect 1285 2421 1319 2455
rect 1149 2335 1183 2369
rect 1217 2335 1251 2369
rect 1285 2335 1319 2369
rect 1149 2249 1183 2283
rect 1217 2249 1251 2283
rect 1285 2249 1319 2283
<< mvndiffc >>
rect 148 2149 182 2183
rect 216 2149 250 2183
rect 284 2149 318 2183
rect 352 2149 386 2183
rect 1149 2054 1183 2088
rect 1217 2054 1251 2088
rect 1285 2054 1319 2088
rect 148 1993 182 2027
rect 216 1993 250 2027
rect 284 1993 318 2027
rect 352 1993 386 2027
rect 148 1837 182 1871
rect 216 1837 250 1871
rect 284 1837 318 1871
rect 352 1837 386 1871
rect 1149 1818 1183 1852
rect 1217 1818 1251 1852
rect 1285 1818 1319 1852
rect 1149 1582 1183 1616
rect 1217 1582 1251 1616
rect 1285 1582 1319 1616
rect 1143 1461 1177 1495
rect 1211 1461 1245 1495
rect 1279 1461 1313 1495
rect 1143 1225 1177 1259
rect 1211 1225 1245 1259
rect 1279 1225 1313 1259
rect 1143 989 1177 1023
rect 1211 989 1245 1023
rect 1279 989 1313 1023
rect 1144 793 1178 827
rect 1212 793 1246 827
rect 1280 793 1314 827
rect 1348 793 1382 827
rect 1144 637 1178 671
rect 1212 637 1246 671
rect 1280 637 1314 671
rect 1348 637 1382 671
rect 1144 481 1178 515
rect 1212 481 1246 515
rect 1280 481 1314 515
rect 1348 481 1382 515
rect 1144 356 1178 390
rect 1212 356 1246 390
rect 1280 356 1314 390
rect 1348 356 1382 390
rect 1144 200 1178 234
rect 1212 200 1246 234
rect 1280 200 1314 234
rect 1348 200 1382 234
rect 1144 44 1178 78
rect 1212 44 1246 78
rect 1280 44 1314 78
rect 1348 44 1382 78
<< mvpdiffc >>
rect 4379 -62 4413 -28
rect 4379 -130 4413 -96
rect 4555 -62 4589 -28
rect 4555 -130 4589 -96
rect 4731 -62 4765 -28
rect 4731 -130 4765 -96
<< psubdiff >>
rect 1530 2073 1564 2097
rect 1530 2005 1564 2039
rect 1530 1937 1564 1971
rect 1530 1869 1564 1903
rect 1530 1801 1564 1835
rect 1530 1733 1564 1767
rect 1530 1665 1564 1699
rect 1530 1597 1564 1631
rect 1530 1529 1564 1563
rect 1530 1461 1564 1495
rect 1530 1393 1564 1427
rect 1530 1325 1564 1359
rect 1530 1257 1564 1291
rect 1530 1189 1564 1223
rect 1530 1121 1564 1155
rect 1530 1052 1564 1087
rect 1530 983 1564 1018
rect 1530 914 1564 949
rect 1530 845 1564 880
rect 1530 776 1564 811
rect 1530 707 1564 742
rect 1530 638 1564 673
rect 1530 569 1564 604
rect 1530 500 1564 535
rect 1530 431 1564 466
rect 1530 362 1564 397
rect 1530 293 1564 328
rect 1530 224 1564 259
rect 1530 155 1564 190
rect 1530 86 1564 121
rect 1530 28 1564 52
<< psubdiffcont >>
rect 1530 2039 1564 2073
rect 1530 1971 1564 2005
rect 1530 1903 1564 1937
rect 1530 1835 1564 1869
rect 1530 1767 1564 1801
rect 1530 1699 1564 1733
rect 1530 1631 1564 1665
rect 1530 1563 1564 1597
rect 1530 1495 1564 1529
rect 1530 1427 1564 1461
rect 1530 1359 1564 1393
rect 1530 1291 1564 1325
rect 1530 1223 1564 1257
rect 1530 1155 1564 1189
rect 1530 1087 1564 1121
rect 1530 1018 1564 1052
rect 1530 949 1564 983
rect 1530 880 1564 914
rect 1530 811 1564 845
rect 1530 742 1564 776
rect 1530 673 1564 707
rect 1530 604 1564 638
rect 1530 535 1564 569
rect 1530 466 1564 500
rect 1530 397 1564 431
rect 1530 328 1564 362
rect 1530 259 1564 293
rect 1530 190 1564 224
rect 1530 121 1564 155
rect 1530 52 1564 86
<< poly >>
rect 1033 2584 1099 2600
rect 1033 2550 1049 2584
rect 1083 2582 1099 2584
rect 1083 2552 1131 2582
rect 1331 2552 1363 2582
rect 1083 2550 1099 2552
rect 1033 2516 1099 2550
rect 1033 2482 1049 2516
rect 1083 2496 1099 2516
rect 1083 2482 1131 2496
rect 1033 2466 1131 2482
rect 1331 2466 1363 2496
rect 1033 2394 1131 2410
rect 1033 2360 1049 2394
rect 1083 2380 1131 2394
rect 1331 2380 1363 2410
rect 1083 2360 1099 2380
rect 1033 2326 1099 2360
rect 1033 2292 1049 2326
rect 1083 2324 1099 2326
rect 1083 2294 1131 2324
rect 1331 2294 1363 2324
rect 1083 2292 1099 2294
rect 1033 2276 1099 2292
rect 0 2122 98 2138
rect 0 2088 16 2122
rect 50 2088 98 2122
rect 0 2038 98 2088
rect 398 2038 430 2138
rect 0 2027 66 2038
rect 0 1993 16 2027
rect 50 1993 66 2027
rect 0 1982 66 1993
rect 1033 2027 1131 2043
rect 1033 1993 1049 2027
rect 1083 1993 1131 2027
rect 0 1932 98 1982
rect 0 1898 16 1932
rect 50 1898 98 1932
rect 0 1882 98 1898
rect 398 1882 430 1982
rect 1033 1954 1131 1993
rect 1033 1920 1049 1954
rect 1083 1920 1131 1954
rect 1033 1881 1131 1920
rect 1033 1847 1049 1881
rect 1083 1863 1131 1881
rect 1331 1863 1363 2043
rect 1083 1847 1099 1863
rect 1033 1808 1099 1847
rect 1033 1774 1049 1808
rect 1083 1807 1099 1808
rect 1083 1774 1131 1807
rect 1033 1735 1131 1774
rect 1033 1701 1049 1735
rect 1083 1701 1131 1735
rect 1033 1662 1131 1701
rect 1033 1628 1049 1662
rect 1083 1628 1131 1662
rect 1033 1627 1131 1628
rect 1331 1627 1363 1807
rect 1033 1589 1099 1627
rect 1033 1555 1049 1589
rect 1083 1555 1099 1589
rect 1033 1516 1099 1555
rect 1033 1482 1049 1516
rect 1083 1482 1099 1516
rect 1033 1450 1099 1482
rect 1033 1444 1131 1450
rect 1033 1410 1049 1444
rect 1083 1410 1131 1444
rect 1033 1372 1131 1410
rect 1033 1338 1049 1372
rect 1083 1338 1131 1372
rect 1033 1300 1131 1338
rect 1033 1266 1049 1300
rect 1083 1270 1131 1300
rect 1331 1270 1363 1450
rect 1083 1266 1099 1270
rect 1033 1228 1099 1266
rect 1033 1194 1049 1228
rect 1083 1214 1099 1228
rect 1083 1194 1131 1214
rect 1033 1156 1131 1194
rect 1033 1122 1049 1156
rect 1083 1122 1131 1156
rect 1033 1084 1131 1122
rect 1033 1050 1049 1084
rect 1083 1050 1131 1084
rect 1033 1034 1131 1050
rect 1331 1034 1363 1214
rect 1034 766 1132 782
rect 1034 732 1050 766
rect 1084 732 1132 766
rect 1034 682 1132 732
rect 1432 682 1464 782
rect 1034 671 1100 682
rect 1034 637 1050 671
rect 1084 637 1100 671
rect 1034 626 1100 637
rect 1034 576 1132 626
rect 1034 542 1050 576
rect 1084 542 1132 576
rect 1034 526 1132 542
rect 1432 526 1464 626
rect 1034 329 1132 345
rect 1034 295 1050 329
rect 1084 295 1132 329
rect 1034 245 1132 295
rect 1432 245 1464 345
rect 1034 234 1100 245
rect 1034 200 1050 234
rect 1084 200 1100 234
rect 1034 189 1100 200
rect 1034 139 1132 189
rect 1034 105 1050 139
rect 1084 105 1132 139
rect 1034 89 1132 105
rect 1432 89 1464 189
rect 4408 80 4544 96
rect 4408 46 4424 80
rect 4458 46 4494 80
rect 4528 46 4544 80
rect 4408 30 4544 46
rect 4424 -2 4544 30
rect 4600 80 4736 96
rect 4600 46 4616 80
rect 4650 46 4686 80
rect 4720 46 4736 80
rect 4600 30 4736 46
rect 4600 -2 4720 30
rect 4424 -174 4544 -142
rect 4600 -174 4720 -142
<< polycont >>
rect 1049 2550 1083 2584
rect 1049 2482 1083 2516
rect 1049 2360 1083 2394
rect 1049 2292 1083 2326
rect 16 2088 50 2122
rect 16 1993 50 2027
rect 1049 1993 1083 2027
rect 16 1898 50 1932
rect 1049 1920 1083 1954
rect 1049 1847 1083 1881
rect 1049 1774 1083 1808
rect 1049 1701 1083 1735
rect 1049 1628 1083 1662
rect 1049 1555 1083 1589
rect 1049 1482 1083 1516
rect 1049 1410 1083 1444
rect 1049 1338 1083 1372
rect 1049 1266 1083 1300
rect 1049 1194 1083 1228
rect 1049 1122 1083 1156
rect 1049 1050 1083 1084
rect 1050 732 1084 766
rect 1050 637 1084 671
rect 1050 542 1084 576
rect 1050 295 1084 329
rect 1050 200 1084 234
rect 1050 105 1084 139
rect 4424 46 4458 80
rect 4494 46 4528 80
rect 4616 46 4650 80
rect 4686 46 4720 80
<< locali >>
rect 1132 2627 1553 2651
rect 1049 2588 1083 2600
rect 1132 2594 1149 2627
rect 1133 2593 1149 2594
rect 1183 2593 1217 2627
rect 1251 2593 1285 2627
rect 1319 2594 1553 2627
rect 1319 2593 1335 2594
rect 1049 2516 1083 2550
rect 1133 2507 1149 2541
rect 1183 2507 1217 2541
rect 1257 2507 1285 2541
rect 1329 2507 1335 2541
rect 1049 2466 1083 2478
rect 1443 2470 1553 2594
rect 1132 2455 1553 2470
rect 1132 2421 1149 2455
rect 1183 2421 1217 2455
rect 1251 2421 1285 2455
rect 1319 2421 1553 2455
rect 1132 2413 1553 2421
rect 1049 2398 1083 2410
rect 1049 2326 1083 2360
rect 1165 2369 1203 2372
rect 1183 2338 1203 2369
rect 1133 2335 1149 2338
rect 1183 2335 1217 2338
rect 1251 2335 1285 2369
rect 1319 2335 1335 2369
rect 132 2183 523 2294
rect 1443 2294 1553 2413
rect 1049 2276 1083 2288
rect 1132 2283 1553 2294
rect 1132 2249 1149 2283
rect 1183 2249 1217 2283
rect 1251 2249 1285 2283
rect 1319 2249 1553 2283
rect 1132 2237 1553 2249
rect 132 2149 148 2183
rect 182 2149 216 2183
rect 250 2149 284 2183
rect 318 2149 352 2183
rect 386 2149 523 2183
rect 132 2148 523 2149
rect 16 2126 50 2138
rect 16 2027 50 2088
rect 1133 2054 1149 2088
rect 1183 2054 1217 2088
rect 1251 2054 1285 2088
rect 1319 2054 1335 2088
rect 1530 2073 1564 2097
rect 1217 2048 1251 2054
rect 1049 2031 1083 2043
rect 298 2027 336 2028
rect 132 1993 148 2027
rect 182 1993 216 2027
rect 250 1994 264 2027
rect 318 1994 336 2027
rect 250 1993 284 1994
rect 318 1993 352 1994
rect 386 1993 402 2027
rect 16 1932 50 1993
rect 16 1882 50 1894
rect 1049 1958 1083 1993
rect 1049 1885 1083 1920
rect 1530 2005 1564 2039
rect 1530 1937 1564 1971
rect 132 1837 148 1871
rect 182 1837 216 1871
rect 250 1837 284 1871
rect 318 1837 352 1871
rect 386 1837 503 1871
rect 134 1702 503 1837
rect 1049 1812 1083 1847
rect 1530 1869 1564 1903
rect 1125 1818 1149 1852
rect 1183 1818 1217 1852
rect 1251 1818 1285 1852
rect 1319 1818 1335 1852
rect 1125 1814 1159 1818
rect 1530 1813 1564 1835
rect 1049 1739 1083 1774
rect 1049 1666 1083 1701
rect 1530 1741 1564 1767
rect 1049 1593 1083 1628
rect 1217 1616 1251 1636
rect 1530 1669 1564 1699
rect 1133 1582 1149 1616
rect 1183 1582 1217 1616
rect 1251 1582 1285 1616
rect 1319 1582 1335 1616
rect 1530 1597 1564 1631
rect 1049 1520 1083 1555
rect 1530 1529 1564 1563
rect 1049 1447 1083 1482
rect 1125 1461 1143 1486
rect 1177 1461 1211 1495
rect 1245 1461 1279 1495
rect 1313 1461 1329 1495
rect 1530 1461 1564 1491
rect 1125 1448 1159 1461
rect 1049 1374 1083 1410
rect 1049 1301 1083 1338
rect 1530 1393 1564 1419
rect 1530 1325 1564 1347
rect 1049 1228 1083 1266
rect 1299 1259 1333 1260
rect 1127 1225 1143 1259
rect 1177 1225 1211 1259
rect 1245 1225 1279 1259
rect 1313 1225 1333 1259
rect 1049 1156 1083 1194
rect 1299 1222 1333 1225
rect 1530 1257 1564 1275
rect 1530 1189 1564 1203
rect 1049 1084 1083 1120
rect 1530 1121 1564 1131
rect 1049 1034 1083 1046
rect 1125 1023 1159 1025
rect 1530 1052 1564 1059
rect 1125 989 1143 1023
rect 1177 989 1211 1023
rect 1245 989 1279 1023
rect 1313 989 1329 1023
rect 1125 987 1159 989
rect 1530 983 1564 987
rect 1530 914 1564 915
rect 1530 877 1564 880
rect 1377 827 1411 828
rect 1128 793 1144 827
rect 1178 793 1212 827
rect 1246 793 1280 827
rect 1314 793 1348 827
rect 1382 793 1411 827
rect 1377 790 1411 793
rect 1050 770 1084 782
rect 1078 766 1084 770
rect 1530 804 1564 811
rect 1044 732 1050 736
rect 1044 671 1084 732
rect 1530 731 1564 742
rect 1218 671 1252 673
rect 1128 637 1144 671
rect 1178 637 1212 671
rect 1246 637 1280 671
rect 1314 637 1348 671
rect 1382 637 1398 671
rect 1530 658 1564 673
rect 1044 576 1084 637
rect 1218 635 1252 637
rect 1044 572 1050 576
rect 1530 585 1564 604
rect 1078 538 1084 542
rect 1050 526 1084 538
rect 1377 515 1411 517
rect 1128 481 1144 515
rect 1178 481 1212 515
rect 1246 481 1280 515
rect 1314 481 1348 515
rect 1382 481 1411 515
rect 1377 479 1411 481
rect 1530 512 1564 535
rect 1530 439 1564 466
rect 1217 390 1251 394
rect 1128 356 1144 390
rect 1178 356 1212 390
rect 1246 356 1280 390
rect 1314 356 1348 390
rect 1382 356 1398 390
rect 1530 366 1564 397
rect 1050 334 1084 345
rect 1077 329 1084 334
rect 1043 295 1050 300
rect 1043 235 1084 295
rect 1530 293 1564 328
rect 1077 234 1084 235
rect 1043 200 1050 201
rect 1043 139 1084 200
rect 1125 234 1159 236
rect 1125 200 1144 234
rect 1178 200 1212 234
rect 1246 200 1280 234
rect 1314 200 1348 234
rect 1382 200 1398 234
rect 1530 224 1564 259
rect 1125 198 1159 200
rect 1043 136 1050 139
rect 1530 155 1564 186
rect 1077 102 1084 105
rect 1050 89 1084 102
rect 1217 78 1251 81
rect 1530 86 1564 113
rect 1128 44 1144 78
rect 1178 44 1212 78
rect 1246 44 1280 78
rect 1314 44 1348 78
rect 1382 44 1398 78
rect 1217 43 1251 44
rect 4408 46 4424 80
rect 4458 46 4494 80
rect 4528 46 4544 80
rect 4600 46 4616 80
rect 4671 62 4686 80
rect 4650 46 4686 62
rect 4720 46 4736 80
rect 1530 28 1564 40
rect 4379 -28 4391 -12
rect 4413 -62 4425 -31
rect 4379 -96 4425 -62
rect 4413 -100 4425 -96
rect 4379 -134 4391 -130
rect 4459 -66 4519 46
rect 4637 24 4671 46
rect 4459 -100 4465 -66
rect 4499 -100 4519 -66
rect 4379 -146 4413 -134
rect 4459 -138 4519 -100
rect 4459 -172 4465 -138
rect 4499 -172 4519 -138
rect 4555 -28 4589 -12
rect 4555 -96 4589 -62
rect 4555 -146 4589 -130
rect 4731 -21 4765 -12
rect 4731 -93 4765 -62
rect 4731 -146 4765 -130
<< viali >>
rect 1049 2584 1083 2588
rect 1049 2554 1083 2584
rect 1049 2482 1083 2512
rect 1223 2507 1251 2541
rect 1251 2507 1257 2541
rect 1295 2507 1319 2541
rect 1319 2507 1329 2541
rect 1049 2478 1083 2482
rect 1049 2394 1083 2398
rect 1049 2364 1083 2394
rect 1131 2369 1165 2372
rect 1203 2369 1237 2372
rect 1131 2338 1149 2369
rect 1149 2338 1165 2369
rect 1203 2338 1217 2369
rect 1217 2338 1237 2369
rect 1049 2292 1083 2322
rect 1049 2288 1083 2292
rect 16 2122 50 2126
rect 16 2092 50 2122
rect 1217 2088 1251 2120
rect 1217 2086 1251 2088
rect 264 2027 298 2028
rect 336 2027 370 2028
rect 1049 2027 1083 2031
rect 16 1993 50 2027
rect 264 1994 284 2027
rect 284 1994 298 2027
rect 336 1994 352 2027
rect 352 1994 370 2027
rect 1049 1997 1083 2027
rect 1217 2014 1251 2048
rect 16 1898 50 1928
rect 16 1894 50 1898
rect 1049 1954 1083 1958
rect 1049 1924 1083 1954
rect 1049 1881 1083 1885
rect 1049 1851 1083 1881
rect 1049 1808 1083 1812
rect 1049 1778 1083 1808
rect 1125 1852 1159 1886
rect 1125 1780 1159 1814
rect 1530 1801 1564 1813
rect 1049 1735 1083 1739
rect 1049 1705 1083 1735
rect 1530 1779 1564 1801
rect 1530 1733 1564 1741
rect 1530 1707 1564 1733
rect 1049 1662 1083 1666
rect 1049 1632 1083 1662
rect 1217 1636 1251 1670
rect 1530 1665 1564 1669
rect 1530 1635 1564 1665
rect 1049 1589 1083 1593
rect 1049 1559 1083 1589
rect 1217 1582 1251 1598
rect 1217 1564 1251 1582
rect 1530 1563 1564 1597
rect 1049 1516 1083 1520
rect 1049 1486 1083 1516
rect 1049 1444 1083 1447
rect 1049 1413 1083 1444
rect 1125 1495 1159 1520
rect 1530 1495 1564 1525
rect 1125 1486 1143 1495
rect 1143 1486 1159 1495
rect 1530 1491 1564 1495
rect 1125 1414 1159 1448
rect 1530 1427 1564 1453
rect 1530 1419 1564 1427
rect 1049 1372 1083 1374
rect 1049 1340 1083 1372
rect 1049 1300 1083 1301
rect 1049 1267 1083 1300
rect 1530 1359 1564 1381
rect 1530 1347 1564 1359
rect 1299 1260 1333 1294
rect 1049 1194 1083 1228
rect 1299 1188 1333 1222
rect 1530 1291 1564 1309
rect 1530 1275 1564 1291
rect 1530 1223 1564 1237
rect 1530 1203 1564 1223
rect 1049 1122 1083 1154
rect 1049 1120 1083 1122
rect 1049 1050 1083 1080
rect 1530 1155 1564 1165
rect 1530 1131 1564 1155
rect 1530 1087 1564 1093
rect 1530 1059 1564 1087
rect 1049 1046 1083 1050
rect 1125 1025 1159 1059
rect 1530 1018 1564 1021
rect 1125 953 1159 987
rect 1530 987 1564 1018
rect 1530 915 1564 949
rect 1377 828 1411 862
rect 1044 766 1078 770
rect 1044 736 1050 766
rect 1050 736 1078 766
rect 1377 756 1411 790
rect 1530 845 1564 877
rect 1530 843 1564 845
rect 1530 776 1564 804
rect 1530 770 1564 776
rect 1530 707 1564 731
rect 1218 673 1252 707
rect 1530 697 1564 707
rect 1044 637 1050 671
rect 1050 637 1078 671
rect 1530 638 1564 658
rect 1218 601 1252 635
rect 1530 624 1564 638
rect 1044 542 1050 572
rect 1050 542 1078 572
rect 1530 569 1564 585
rect 1530 551 1564 569
rect 1044 538 1078 542
rect 1377 517 1411 551
rect 1377 445 1411 479
rect 1530 500 1564 512
rect 1530 478 1564 500
rect 1530 431 1564 439
rect 1217 394 1251 428
rect 1530 405 1564 431
rect 1530 362 1564 366
rect 1043 329 1077 334
rect 1043 300 1050 329
rect 1050 300 1077 329
rect 1217 322 1251 356
rect 1530 332 1564 362
rect 1043 234 1077 235
rect 1043 201 1050 234
rect 1050 201 1077 234
rect 1125 236 1159 270
rect 1530 259 1564 293
rect 1125 164 1159 198
rect 1530 190 1564 220
rect 1530 186 1564 190
rect 1043 105 1050 136
rect 1050 105 1077 136
rect 1530 121 1564 147
rect 1043 102 1077 105
rect 1217 81 1251 115
rect 1530 113 1564 121
rect 4637 80 4671 96
rect 1530 52 1564 74
rect 1217 9 1251 43
rect 1530 40 1564 52
rect 4637 62 4650 80
rect 4650 62 4671 80
rect 4391 -28 4425 3
rect 4391 -31 4413 -28
rect 4413 -31 4425 -28
rect 4391 -130 4413 -100
rect 4413 -130 4425 -100
rect 4391 -134 4425 -130
rect 4637 -10 4671 24
rect 4465 -100 4499 -66
rect 4465 -172 4499 -138
rect 4731 -28 4765 -21
rect 4731 -55 4765 -28
rect 4731 -96 4765 -93
rect 4731 -127 4765 -96
<< metal1 >>
rect 1043 2588 1089 2600
rect 1043 2554 1049 2588
rect 1083 2554 1089 2588
rect 1043 2512 1089 2554
rect 1043 2478 1049 2512
rect 1083 2478 1089 2512
rect 1211 2541 1341 2547
rect 1211 2507 1223 2541
rect 1257 2507 1295 2541
rect 1329 2507 1341 2541
rect 1211 2501 1341 2507
rect 1043 2466 1089 2478
rect 1043 2398 1089 2410
rect 1043 2364 1049 2398
rect 1083 2364 1089 2398
rect 1043 2322 1089 2364
rect 1043 2288 1049 2322
rect 1083 2288 1089 2322
rect 1043 2276 1089 2288
rect 1119 2372 1249 2378
rect 1119 2338 1131 2372
rect 1165 2338 1203 2372
rect 1237 2338 1249 2372
rect 1119 2332 1249 2338
rect 10 2126 56 2138
rect 10 2092 16 2126
rect 50 2092 56 2126
rect 10 2027 56 2092
rect 10 1993 16 2027
rect 50 1993 56 2027
rect 10 1928 56 1993
rect 251 1985 257 2037
rect 309 1985 324 2037
rect 376 1985 382 2037
rect 1043 2031 1089 2043
rect 1043 1997 1049 2031
rect 1083 1997 1089 2031
rect 10 1894 16 1928
rect 50 1894 56 1928
rect 10 1882 56 1894
rect 1043 1958 1089 1997
rect 1043 1924 1049 1958
rect 1083 1924 1089 1958
rect 1043 1885 1089 1924
rect 1043 1851 1049 1885
rect 1083 1851 1089 1885
rect 1043 1812 1089 1851
rect 1043 1778 1049 1812
rect 1083 1778 1089 1812
rect 1043 1739 1089 1778
rect 1119 1886 1165 2332
rect 1119 1852 1125 1886
rect 1159 1852 1165 1886
rect 1119 1814 1165 1852
rect 1119 1780 1125 1814
rect 1159 1780 1165 1814
rect 1119 1768 1165 1780
rect 1211 2120 1257 2132
rect 1211 2086 1217 2120
rect 1251 2086 1257 2120
rect 1211 2048 1257 2086
rect 1211 2014 1217 2048
rect 1251 2014 1257 2048
rect 1043 1705 1049 1739
rect 1083 1705 1089 1739
rect 1043 1666 1089 1705
rect 1043 1632 1049 1666
rect 1083 1632 1089 1666
rect 1043 1593 1089 1632
rect 1043 1559 1049 1593
rect 1083 1559 1089 1593
rect 1043 1520 1089 1559
rect 1211 1670 1257 2014
rect 1211 1636 1217 1670
rect 1251 1636 1257 1670
rect 1211 1598 1257 1636
rect 1211 1564 1217 1598
rect 1251 1564 1257 1598
rect 1043 1486 1049 1520
rect 1083 1486 1089 1520
rect 1043 1447 1089 1486
rect 1043 1413 1049 1447
rect 1083 1413 1089 1447
rect 1043 1374 1089 1413
rect 1043 1340 1049 1374
rect 1083 1340 1089 1374
rect 1043 1301 1089 1340
rect 1043 1267 1049 1301
rect 1083 1267 1089 1301
rect 1043 1228 1089 1267
rect 1043 1194 1049 1228
rect 1083 1194 1089 1228
rect 1043 1154 1089 1194
rect 1043 1120 1049 1154
rect 1083 1120 1089 1154
rect 1043 1080 1089 1120
rect 1043 1046 1049 1080
rect 1083 1046 1089 1080
rect 1043 1034 1089 1046
rect 1119 1520 1165 1532
rect 1119 1486 1125 1520
rect 1159 1486 1165 1520
rect 1119 1448 1165 1486
rect 1119 1414 1125 1448
rect 1159 1414 1165 1448
rect 1119 1059 1165 1414
rect 1119 1025 1125 1059
rect 1159 1025 1165 1059
rect 1119 987 1165 1025
rect 1119 953 1125 987
rect 1159 953 1165 987
rect 1038 770 1084 782
rect 1038 736 1044 770
rect 1078 736 1084 770
rect 1038 671 1084 736
rect 1038 637 1044 671
rect 1078 637 1084 671
rect 1038 572 1084 637
rect 1038 538 1044 572
rect 1078 538 1084 572
rect 1038 526 1084 538
rect 1037 334 1083 526
rect 1037 300 1043 334
rect 1077 300 1083 334
rect 1037 235 1083 300
rect 1037 201 1043 235
rect 1077 201 1083 235
rect 1037 136 1083 201
rect 1119 270 1165 953
rect 1211 719 1257 1564
rect 1293 1294 1339 2501
rect 1293 1260 1299 1294
rect 1333 1260 1339 1294
rect 1293 1222 1339 1260
rect 1293 1188 1299 1222
rect 1333 1188 1339 1222
rect 1293 1176 1339 1188
rect 1371 1985 1377 2037
rect 1429 1985 1441 2037
rect 1493 1985 1499 2037
rect 1371 862 1417 1985
rect 1371 828 1377 862
rect 1411 828 1417 862
rect 1371 790 1417 828
rect 1371 756 1377 790
rect 1411 756 1417 790
rect 1211 707 1258 719
rect 1211 673 1218 707
rect 1252 673 1258 707
rect 1211 645 1258 673
rect 1212 635 1258 645
rect 1212 601 1218 635
rect 1252 601 1258 635
rect 1212 589 1258 601
rect 1371 551 1417 756
rect 1371 535 1377 551
rect 1411 535 1417 551
rect 1524 1813 1570 1825
rect 1524 1779 1530 1813
rect 1564 1779 1570 1813
rect 1524 1741 1570 1779
rect 1524 1707 1530 1741
rect 1564 1707 1570 1741
rect 1524 1669 1570 1707
rect 1524 1635 1530 1669
rect 1564 1635 1570 1669
rect 1524 1597 1570 1635
rect 1524 1563 1530 1597
rect 1564 1563 1570 1597
rect 1524 1525 1570 1563
rect 1524 1491 1530 1525
rect 1564 1491 1570 1525
rect 1524 1453 1570 1491
rect 1524 1419 1530 1453
rect 1564 1419 1570 1453
rect 1524 1381 1570 1419
rect 1524 1347 1530 1381
rect 1564 1347 1570 1381
rect 1524 1309 1570 1347
rect 1524 1275 1530 1309
rect 1564 1275 1570 1309
rect 1524 1237 1570 1275
rect 1524 1203 1530 1237
rect 1564 1203 1570 1237
rect 1524 1165 1570 1203
rect 1524 1131 1530 1165
rect 1564 1131 1570 1165
rect 1524 1093 1570 1131
rect 1524 1059 1530 1093
rect 1564 1059 1570 1093
rect 1524 1021 1570 1059
rect 1524 987 1530 1021
rect 1564 987 1570 1021
rect 1524 949 1570 987
rect 1524 915 1530 949
rect 1564 915 1570 949
rect 1524 877 1570 915
rect 1524 843 1530 877
rect 1564 843 1570 877
rect 1524 804 1570 843
rect 1524 770 1530 804
rect 1564 770 1570 804
rect 1524 731 1570 770
rect 1524 697 1530 731
rect 1564 697 1570 731
rect 1524 658 1570 697
rect 1524 624 1530 658
rect 1564 624 1570 658
rect 1524 585 1570 624
rect 1524 551 1530 585
rect 1564 551 1570 585
rect 4568 567 4574 619
rect 4626 567 4638 619
rect 4690 567 4696 619
rect 1293 483 1299 535
rect 1351 483 1363 535
rect 1415 483 1421 535
rect 1524 512 1570 551
rect 1371 479 1417 483
rect 1203 394 1209 446
rect 1261 394 1273 446
rect 1325 394 1331 446
rect 1371 445 1377 479
rect 1411 445 1417 479
rect 1371 433 1417 445
rect 1524 478 1530 512
rect 1564 478 1570 512
rect 1524 439 1570 478
rect 1524 405 1530 439
rect 1564 405 1570 439
rect 1119 236 1125 270
rect 1159 236 1165 270
rect 1119 198 1165 236
rect 1119 164 1125 198
rect 1159 164 1165 198
rect 1119 152 1165 164
rect 1211 356 1257 394
rect 1211 322 1217 356
rect 1251 322 1257 356
rect 1037 102 1043 136
rect 1077 102 1083 136
rect 1037 90 1083 102
rect 1211 115 1257 322
rect 1211 81 1217 115
rect 1251 81 1257 115
rect 1211 43 1257 81
rect 1211 9 1217 43
rect 1251 9 1257 43
rect 1524 366 1570 405
rect 1524 332 1530 366
rect 1564 332 1570 366
rect 1524 293 1570 332
rect 1524 259 1530 293
rect 1564 259 1570 293
rect 1524 220 1570 259
rect 1524 186 1530 220
rect 1564 186 1570 220
rect 1524 147 1570 186
rect 1524 113 1530 147
rect 1564 113 1570 147
rect 1524 74 1570 113
rect 4663 108 4696 567
rect 1524 40 1530 74
rect 1564 40 1570 74
rect 4631 96 4696 108
rect 4631 62 4637 96
rect 4671 62 4696 96
rect 1524 28 1570 40
tri 4614 28 4631 45 se
rect 4631 28 4696 62
tri 4610 24 4614 28 se
rect 4614 24 4696 28
tri 4601 15 4610 24 se
rect 4610 15 4637 24
rect 1211 -3 1257 9
rect 4385 3 4637 15
rect 4385 -31 4391 3
rect 4425 -10 4637 3
rect 4671 -10 4696 24
rect 4860 600 4912 606
rect 4860 536 4912 548
rect 4860 403 4912 484
rect 4425 -22 4696 -10
rect 4725 -21 4771 -9
rect 4425 -31 4431 -22
rect 4385 -100 4431 -31
tri 4431 -39 4448 -22 nw
rect 4725 -54 4731 -21
rect 4385 -134 4391 -100
rect 4425 -134 4431 -100
rect 4385 -146 4431 -134
rect 4459 -55 4731 -54
rect 4765 -54 4771 -21
tri 4857 -22 4860 -19 se
rect 4860 -22 4893 403
tri 4893 384 4912 403 nw
tri 4825 -54 4857 -22 se
rect 4857 -54 4893 -22
rect 4765 -55 4893 -54
rect 4459 -66 4893 -55
rect 4459 -100 4465 -66
rect 4499 -93 4893 -66
rect 4499 -100 4731 -93
rect 4459 -127 4731 -100
rect 4765 -127 4893 -93
rect 4459 -133 4893 -127
rect 4459 -138 4505 -133
rect 4459 -172 4465 -138
rect 4499 -172 4505 -138
rect 4725 -139 4771 -133
tri 4828 -139 4834 -133 ne
rect 4834 -139 4893 -133
tri 4834 -166 4861 -139 ne
rect 4861 -165 4893 -139
rect 4459 -184 4505 -172
<< via1 >>
rect 257 2028 309 2037
rect 257 1994 264 2028
rect 264 1994 298 2028
rect 298 1994 309 2028
rect 257 1985 309 1994
rect 324 2028 376 2037
rect 324 1994 336 2028
rect 336 1994 370 2028
rect 370 1994 376 2028
rect 324 1985 376 1994
rect 1377 1985 1429 2037
rect 1441 1985 1493 2037
rect 4574 567 4626 619
rect 4638 567 4690 619
rect 1299 483 1351 535
rect 1363 517 1377 535
rect 1377 517 1411 535
rect 1411 517 1415 535
rect 1363 483 1415 517
rect 1209 428 1261 446
rect 1209 394 1217 428
rect 1217 394 1251 428
rect 1251 394 1261 428
rect 1273 394 1325 446
rect 4860 548 4912 600
rect 4860 484 4912 536
<< metal2 >>
rect 251 1985 257 2037
rect 309 1985 324 2037
rect 376 1985 1377 2037
rect 1429 1985 1441 2037
rect 1493 1985 1499 2037
tri 4145 567 4197 619 se
rect 4197 567 4574 619
rect 4626 567 4638 619
rect 4690 567 4696 619
rect 4860 600 4912 606
tri 4126 548 4145 567 se
rect 4145 548 4221 567
tri 4221 548 4240 567 nw
tri 4114 536 4126 548 se
rect 4126 536 4209 548
tri 4209 536 4221 548 nw
rect 4860 536 4912 548
tri 4113 535 4114 536 se
rect 4114 535 4208 536
tri 4208 535 4209 536 nw
rect 1293 483 1299 535
rect 1351 483 1363 535
rect 1415 530 4203 535
tri 4203 530 4208 535 nw
rect 1415 529 4202 530
tri 4202 529 4203 530 nw
tri 4285 529 4286 530 se
rect 4286 529 4860 530
rect 1415 484 4157 529
tri 4157 484 4202 529 nw
tri 4240 484 4285 529 se
rect 4285 484 4860 529
rect 1415 483 4156 484
tri 4156 483 4157 484 nw
tri 4239 483 4240 484 se
rect 4240 483 4912 484
tri 4202 446 4239 483 se
rect 4239 478 4912 483
rect 4239 446 4297 478
tri 4297 446 4329 478 nw
rect 1203 394 1209 446
rect 1261 394 1273 446
rect 1325 394 4245 446
tri 4245 394 4297 446 nw
use sky130_fd_pr__nfet_01v8__example_55959141808496  sky130_fd_pr__nfet_01v8__example_55959141808496_0
timestamp 1663361622
transform 0 1 1131 1 0 1034
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808497  sky130_fd_pr__nfet_01v8__example_55959141808497_0
timestamp 1663361622
transform 0 -1 1331 1 0 1627
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808502  sky130_fd_pr__nfet_01v8__example_55959141808502_0
timestamp 1663361622
transform 0 -1 1331 1 0 2294
box -1 0 289 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_0
timestamp 1663361622
transform 0 1 1132 1 0 526
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_1
timestamp 1663361622
transform 0 1 1132 1 0 89
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_2
timestamp 1663361622
transform 0 -1 398 -1 0 2138
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808500  sky130_fd_pr__pfet_01v8__example_55959141808500_0
timestamp 1663361622
transform 1 0 4424 0 1 -142
box -1 0 297 1
<< labels >>
flabel comment s 1060 2348 1060 2348 0 FreeSans 400 90 0 0 IN_H
<< properties >>
string GDS_END 29655542
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 29636978
<< end >>
