magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 1 2 1 3 6 DRAIN
port 2 nsew
rlabel  s 0 3 1 4 4 GATE
port 3 nsew
rlabel  s 1 0 1 3 6 SOURCE
port 4 nsew
rlabel  s 0 0 0 3 4 SOURCE
port 4 nsew
rlabel  s 0 0 1 0 2 SOURCE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 1 4
string LEFview TRUE
<< end >>
