magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 211 157 397 203
rect 30 21 397 157
rect 30 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 108 47 138 131
rect 192 47 222 131
rect 289 47 319 177
<< scpmoshvt >>
rect 120 297 150 381
rect 192 297 222 381
rect 289 297 319 497
<< ndiff >>
rect 237 131 289 177
rect 56 103 108 131
rect 56 69 64 103
rect 98 69 108 103
rect 56 47 108 69
rect 138 103 192 131
rect 138 69 148 103
rect 182 69 192 103
rect 138 47 192 69
rect 222 103 289 131
rect 222 69 244 103
rect 278 69 289 103
rect 222 47 289 69
rect 319 163 371 177
rect 319 129 329 163
rect 363 129 371 163
rect 319 95 371 129
rect 319 61 329 95
rect 363 61 371 95
rect 319 47 371 61
<< pdiff >>
rect 237 469 289 497
rect 237 435 245 469
rect 279 435 289 469
rect 237 401 289 435
rect 237 381 245 401
rect 68 349 120 381
rect 68 315 76 349
rect 110 315 120 349
rect 68 297 120 315
rect 150 297 192 381
rect 222 367 245 381
rect 279 367 289 401
rect 222 297 289 367
rect 319 485 387 497
rect 319 451 345 485
rect 379 451 387 485
rect 319 417 387 451
rect 319 383 345 417
rect 379 383 387 417
rect 319 297 387 383
<< ndiffc >>
rect 64 69 98 103
rect 148 69 182 103
rect 244 69 278 103
rect 329 129 363 163
rect 329 61 363 95
<< pdiffc >>
rect 245 435 279 469
rect 76 315 110 349
rect 245 367 279 401
rect 345 451 379 485
rect 345 383 379 417
<< poly >>
rect 289 497 319 523
rect 120 381 150 407
rect 192 381 222 407
rect 120 265 150 297
rect 50 249 150 265
rect 50 215 66 249
rect 100 215 150 249
rect 50 199 150 215
rect 192 265 222 297
rect 289 265 319 297
rect 192 249 246 265
rect 192 215 202 249
rect 236 215 246 249
rect 192 199 246 215
rect 289 249 355 265
rect 289 215 305 249
rect 339 215 355 249
rect 289 199 355 215
rect 108 131 138 199
rect 192 131 222 199
rect 289 177 319 199
rect 108 21 138 47
rect 192 21 222 47
rect 289 21 319 47
<< polycont >>
rect 66 215 100 249
rect 202 215 236 249
rect 305 215 339 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 229 469 295 527
rect 229 435 245 469
rect 279 435 295 469
rect 229 401 295 435
rect 54 349 132 368
rect 229 367 245 401
rect 279 367 295 401
rect 329 485 436 493
rect 329 451 345 485
rect 379 451 436 485
rect 329 417 436 451
rect 329 383 345 417
rect 379 383 436 417
rect 329 369 436 383
rect 54 315 76 349
rect 110 333 132 349
rect 110 315 339 333
rect 54 299 339 315
rect 29 249 100 265
rect 29 215 66 249
rect 29 153 100 215
rect 134 119 168 299
rect 202 249 255 265
rect 236 215 255 249
rect 202 153 255 215
rect 305 249 339 299
rect 305 199 339 215
rect 373 165 436 369
rect 313 163 436 165
rect 313 129 329 163
rect 363 129 436 163
rect 50 103 98 119
rect 50 69 64 103
rect 50 17 98 69
rect 134 103 190 119
rect 134 69 148 103
rect 182 69 190 103
rect 134 53 190 69
rect 236 103 279 119
rect 236 69 244 103
rect 278 69 279 103
rect 236 17 279 69
rect 313 95 436 129
rect 313 61 329 95
rect 363 61 436 95
rect 313 51 436 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 397 357 431 391 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 or2_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 984256
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 980090
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 2.300 0.000 
<< end >>
