/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/cdl/sky130_fd_sc_hvl/sky130_fd_sc_hvl.cdl