/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__npn_05v5_W1p00L2p00.model.spice