magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1169 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
rect 959 47 989 177
rect 1043 47 1073 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 531 297 561 497
rect 615 297 645 497
rect 699 297 729 497
rect 783 297 813 497
rect 975 297 1005 497
rect 1059 297 1089 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 93 79 131
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 47 163 131
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 165 331 177
rect 277 131 287 165
rect 321 131 331 165
rect 277 47 331 131
rect 361 93 415 177
rect 361 59 371 93
rect 405 59 415 93
rect 361 47 415 59
rect 445 93 603 177
rect 445 59 540 93
rect 574 59 603 93
rect 445 47 603 59
rect 633 165 687 177
rect 633 131 643 165
rect 677 131 687 165
rect 633 93 687 131
rect 633 59 643 93
rect 677 59 687 93
rect 633 47 687 59
rect 717 93 771 177
rect 717 59 727 93
rect 761 59 771 93
rect 717 47 771 59
rect 801 165 959 177
rect 801 131 827 165
rect 861 131 895 165
rect 929 131 959 165
rect 801 93 959 131
rect 801 59 827 93
rect 861 59 895 93
rect 929 59 959 93
rect 801 47 959 59
rect 989 93 1043 177
rect 989 59 999 93
rect 1033 59 1043 93
rect 989 47 1043 59
rect 1073 165 1143 177
rect 1073 131 1101 165
rect 1135 131 1143 165
rect 1073 93 1143 131
rect 1073 59 1101 93
rect 1135 59 1143 93
rect 1073 47 1143 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 417 163 497
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 297 331 451
rect 361 485 413 497
rect 361 451 371 485
rect 405 451 413 485
rect 361 417 413 451
rect 361 383 371 417
rect 405 383 413 417
rect 361 297 413 383
rect 475 485 531 497
rect 475 451 483 485
rect 517 451 531 485
rect 475 417 531 451
rect 475 383 483 417
rect 517 383 531 417
rect 475 297 531 383
rect 561 417 615 497
rect 561 383 571 417
rect 605 383 615 417
rect 561 349 615 383
rect 561 315 571 349
rect 605 315 615 349
rect 561 297 615 315
rect 645 485 699 497
rect 645 451 655 485
rect 689 451 699 485
rect 645 417 699 451
rect 645 383 655 417
rect 689 383 699 417
rect 645 349 699 383
rect 645 315 655 349
rect 689 315 699 349
rect 645 297 699 315
rect 729 417 783 497
rect 729 383 739 417
rect 773 383 783 417
rect 729 349 783 383
rect 729 315 739 349
rect 773 315 783 349
rect 729 297 783 315
rect 813 485 869 497
rect 813 451 827 485
rect 861 451 869 485
rect 813 417 869 451
rect 813 383 827 417
rect 861 383 869 417
rect 813 297 869 383
rect 923 485 975 497
rect 923 451 931 485
rect 965 451 975 485
rect 923 417 975 451
rect 923 383 931 417
rect 965 383 975 417
rect 923 297 975 383
rect 1005 485 1059 497
rect 1005 451 1015 485
rect 1049 451 1059 485
rect 1005 417 1059 451
rect 1005 383 1015 417
rect 1049 383 1059 417
rect 1005 349 1059 383
rect 1005 315 1015 349
rect 1049 315 1059 349
rect 1005 297 1059 315
rect 1089 485 1145 497
rect 1089 451 1103 485
rect 1137 451 1145 485
rect 1089 417 1145 451
rect 1089 383 1103 417
rect 1137 383 1145 417
rect 1089 349 1145 383
rect 1089 315 1103 349
rect 1137 315 1145 349
rect 1089 297 1145 315
<< ndiffc >>
rect 35 131 69 165
rect 35 59 69 93
rect 119 131 153 165
rect 203 59 237 93
rect 287 131 321 165
rect 371 59 405 93
rect 540 59 574 93
rect 643 131 677 165
rect 643 59 677 93
rect 727 59 761 93
rect 827 131 861 165
rect 895 131 929 165
rect 827 59 861 93
rect 895 59 929 93
rect 999 59 1033 93
rect 1101 131 1135 165
rect 1101 59 1135 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 371 451 405 485
rect 371 383 405 417
rect 483 451 517 485
rect 483 383 517 417
rect 571 383 605 417
rect 571 315 605 349
rect 655 451 689 485
rect 655 383 689 417
rect 655 315 689 349
rect 739 383 773 417
rect 739 315 773 349
rect 827 451 861 485
rect 827 383 861 417
rect 931 451 965 485
rect 931 383 965 417
rect 1015 451 1049 485
rect 1015 383 1049 417
rect 1015 315 1049 349
rect 1103 451 1137 485
rect 1103 383 1137 417
rect 1103 315 1137 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 531 497 561 523
rect 615 497 645 523
rect 699 497 729 523
rect 783 497 813 523
rect 975 497 1005 523
rect 1059 497 1089 523
rect 79 265 109 297
rect 163 265 193 297
rect 79 249 193 265
rect 79 215 119 249
rect 153 215 193 249
rect 79 199 193 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 265 277 297
rect 331 265 361 297
rect 247 249 361 265
rect 531 265 561 297
rect 615 265 645 297
rect 699 265 729 297
rect 783 265 813 297
rect 975 265 1005 297
rect 1059 265 1089 297
rect 531 253 645 265
rect 247 215 287 249
rect 321 215 361 249
rect 247 199 361 215
rect 247 177 277 199
rect 331 177 361 199
rect 415 249 645 253
rect 415 223 563 249
rect 415 177 445 223
rect 531 215 563 223
rect 597 215 645 249
rect 531 199 645 215
rect 687 249 813 265
rect 687 215 731 249
rect 765 215 813 249
rect 687 199 813 215
rect 959 249 1089 265
rect 959 215 1001 249
rect 1035 215 1089 249
rect 959 199 1089 215
rect 603 177 633 199
rect 687 177 717 199
rect 771 177 801 199
rect 959 177 989 199
rect 1043 177 1073 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
rect 959 21 989 47
rect 1043 21 1073 47
<< polycont >>
rect 119 215 153 249
rect 287 215 321 249
rect 563 215 597 249
rect 731 215 765 249
rect 1001 215 1035 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 485 253 493
rect 18 451 35 485
rect 69 459 203 485
rect 18 417 69 451
rect 237 451 253 485
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 417 169 419
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 417 253 451
rect 287 485 321 527
rect 287 435 321 451
rect 355 485 421 491
rect 355 451 371 485
rect 405 451 421 485
rect 237 401 253 417
rect 355 417 421 451
rect 355 401 371 417
rect 237 383 371 401
rect 405 383 421 417
rect 203 367 421 383
rect 467 485 877 489
rect 467 451 483 485
rect 517 451 655 485
rect 689 451 827 485
rect 861 451 877 485
rect 467 417 517 451
rect 655 417 689 451
rect 827 417 877 451
rect 467 383 483 417
rect 467 367 517 383
rect 555 383 571 417
rect 605 383 621 417
rect 103 315 119 349
rect 153 333 169 349
rect 555 349 621 383
rect 555 333 571 349
rect 153 315 571 333
rect 605 315 621 349
rect 103 299 621 315
rect 655 349 689 383
rect 655 299 689 315
rect 723 383 739 417
rect 773 383 789 417
rect 723 349 789 383
rect 861 383 877 417
rect 827 367 877 383
rect 924 485 965 527
rect 924 451 931 485
rect 924 417 965 451
rect 924 383 931 417
rect 924 367 965 383
rect 999 485 1065 492
rect 999 451 1015 485
rect 1049 451 1065 485
rect 999 417 1065 451
rect 999 383 1015 417
rect 1049 383 1065 417
rect 723 315 739 349
rect 773 333 789 349
rect 999 349 1065 383
rect 999 333 1015 349
rect 773 315 1015 333
rect 1049 315 1065 349
rect 723 299 1065 315
rect 1099 485 1143 527
rect 1099 451 1103 485
rect 1137 451 1143 485
rect 1099 417 1143 451
rect 1099 383 1103 417
rect 1137 383 1143 417
rect 1099 349 1143 383
rect 1099 315 1103 349
rect 1137 315 1143 349
rect 1099 299 1143 315
rect 18 249 169 265
rect 18 215 119 249
rect 153 215 169 249
rect 203 249 341 265
rect 203 215 287 249
rect 321 215 341 249
rect 375 221 434 299
rect 481 249 613 265
rect 375 181 409 221
rect 481 215 563 249
rect 597 215 613 249
rect 674 249 896 265
rect 674 215 731 249
rect 765 215 896 249
rect 950 249 1173 265
rect 950 215 1001 249
rect 1035 215 1173 249
rect 18 165 69 181
rect 18 131 35 165
rect 103 165 409 181
rect 103 131 119 165
rect 153 131 287 165
rect 321 131 409 165
rect 447 165 1151 181
rect 447 143 643 165
rect 18 97 69 131
rect 447 97 481 143
rect 627 131 643 143
rect 677 143 827 165
rect 677 131 693 143
rect 18 93 481 97
rect 18 59 35 93
rect 69 59 203 93
rect 237 59 371 93
rect 405 59 481 93
rect 18 51 481 59
rect 524 93 590 109
rect 524 59 540 93
rect 574 59 590 93
rect 524 17 590 59
rect 627 93 693 131
rect 811 131 827 143
rect 861 131 895 165
rect 929 143 1101 165
rect 929 131 945 143
rect 627 59 643 93
rect 677 59 693 93
rect 627 51 693 59
rect 727 93 761 109
rect 727 17 761 59
rect 811 93 945 131
rect 1085 131 1101 143
rect 1135 131 1151 165
rect 811 59 827 93
rect 861 59 895 93
rect 929 59 945 93
rect 811 51 945 59
rect 981 93 1047 109
rect 981 59 999 93
rect 1033 59 1047 93
rect 981 17 1047 59
rect 1085 93 1151 131
rect 1085 59 1101 93
rect 1135 59 1151 93
rect 1085 51 1151 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1134 221 1168 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 398 289 432 323 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o32ai_2
rlabel metal1 s 0 -48 1196 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 1497588
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1487662
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.980 0.000 
<< end >>
