/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/fixed_devices/sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4_top_fail.cdl