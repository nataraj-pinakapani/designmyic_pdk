magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel rotate s 4 4 4 4 6 BULK
port 1 nsew
rlabel rotate s 4 3 4 3 6 BULK
port 1 nsew
rlabel rotate s 4 3 4 3 6 BULK
port 1 nsew
rlabel rotate s 4 3 4 3 6 BULK
port 1 nsew
rlabel rotate s 4 2 4 2 6 BULK
port 1 nsew
rlabel rotate s 4 2 4 2 6 BULK
port 1 nsew
rlabel rotate s 4 1 4 2 6 BULK
port 1 nsew
rlabel rotate s 4 1 4 1 6 BULK
port 1 nsew
rlabel rotate s 0 4 0 4 4 BULK
port 1 nsew
rlabel rotate s 0 3 0 3 4 BULK
port 1 nsew
rlabel rotate s 0 3 0 3 4 BULK
port 1 nsew
rlabel rotate s 0 3 0 3 4 BULK
port 1 nsew
rlabel rotate s 0 2 0 2 4 BULK
port 1 nsew
rlabel rotate s 0 2 0 2 4 BULK
port 1 nsew
rlabel rotate s 0 1 0 2 4 BULK
port 1 nsew
rlabel rotate s 0 1 0 1 4 BULK
port 1 nsew
rlabel  s 4 4 4 4 6 BULK
port 1 nsew
rlabel  s 4 1 4 4 6 BULK
port 1 nsew
rlabel  s 4 1 4 1 6 BULK
port 1 nsew
rlabel  s 3 4 4 4 6 BULK
port 1 nsew
rlabel  s 3 0 4 1 8 BULK
port 1 nsew
rlabel  s 1 4 1 4 6 BULK
port 1 nsew
rlabel  s 1 4 1 4 6 BULK
port 1 nsew
rlabel  s 1 1 1 1 6 BULK
port 1 nsew
rlabel  s 1 0 1 1 8 BULK
port 1 nsew
rlabel  s 0 1 1 4 4 BULK
port 1 nsew
rlabel  s 4 1 4 4 6 BULK
port 1 nsew
rlabel  s 0 1 1 4 4 BULK
port 1 nsew
rlabel  s 0 3 4 4 6 DRAIN
port 2 nsew
rlabel rotate s 1 4 3 5 6 GATE
port 3 nsew
rlabel rotate s 1 0 3 1 8 GATE
port 3 nsew
rlabel  s 1 4 3 5 6 GATE
port 3 nsew
rlabel  s 1 0 3 1 8 GATE
port 3 nsew
rlabel  s 1 4 3 5 6 GATE
port 3 nsew
rlabel  s 1 0 3 1 8 GATE
port 3 nsew
rlabel  s 0 1 4 2 6 SOURCE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 4 5
string LEFview TRUE
<< end >>
