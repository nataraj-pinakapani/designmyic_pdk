/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.tech/klayout/lvs/testing/testcases/sky130_fd_pr__nfet_g5v0d10v5_fail.cdl