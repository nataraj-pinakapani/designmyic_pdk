magic
tech minimum
timestamp 1644097874
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -3 -3 4 18
string LEFview TRUE
<< end >>
