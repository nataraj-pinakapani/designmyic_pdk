magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 0 1 30 4 D
port 1 nsew
rlabel  s 6 33 6 36 6 PSUB
port 2 nsew
rlabel  s 6 -3 6 -3 8 PSUB
port 2 nsew
rlabel  s 6 -6 6 -3 8 PSUB
port 2 nsew
rlabel  s -6 36 6 36 4 PSUB
port 2 nsew
rlabel  s -6 33 -5 36 4 PSUB
port 2 nsew
rlabel  s -6 -6 -5 -3 2 PSUB
port 2 nsew
rlabel  s -6 -6 6 -6 2 PSUB
port 2 nsew
rlabel  s -5 0 -5 30 4 S
port 3 nsew
rlabel  s 5 0 6 30 6 S
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -6 -6 6 36
string LEFview TRUE
<< end >>
