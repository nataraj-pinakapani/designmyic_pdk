magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 9 67 1195 203
rect 29 -17 63 67
rect 294 21 1195 67
<< scnmos >>
rect 87 93 117 177
rect 171 93 201 177
rect 388 47 418 177
rect 472 47 502 177
rect 556 47 586 177
rect 640 47 670 177
rect 832 47 862 177
rect 916 47 946 177
rect 1000 47 1030 177
rect 1084 47 1114 177
<< scpmoshvt >>
rect 79 410 109 494
rect 176 297 206 381
rect 388 297 418 497
rect 472 297 502 497
rect 556 297 586 497
rect 640 297 670 497
rect 832 297 862 497
rect 916 297 946 497
rect 1000 297 1030 497
rect 1084 297 1114 497
<< ndiff >>
rect 35 149 87 177
rect 35 115 43 149
rect 77 115 87 149
rect 35 93 87 115
rect 117 149 171 177
rect 117 115 127 149
rect 161 115 171 149
rect 117 93 171 115
rect 201 149 253 177
rect 201 115 211 149
rect 245 115 253 149
rect 201 93 253 115
rect 320 95 388 177
rect 320 61 328 95
rect 362 61 388 95
rect 320 47 388 61
rect 418 163 472 177
rect 418 129 428 163
rect 462 129 472 163
rect 418 95 472 129
rect 418 61 428 95
rect 462 61 472 95
rect 418 47 472 61
rect 502 95 556 177
rect 502 61 512 95
rect 546 61 556 95
rect 502 47 556 61
rect 586 163 640 177
rect 586 129 596 163
rect 630 129 640 163
rect 586 95 640 129
rect 586 61 596 95
rect 630 61 640 95
rect 586 47 640 61
rect 670 95 722 177
rect 670 61 680 95
rect 714 61 722 95
rect 670 47 722 61
rect 776 95 832 177
rect 776 61 788 95
rect 822 61 832 95
rect 776 47 832 61
rect 862 163 916 177
rect 862 129 872 163
rect 906 129 916 163
rect 862 95 916 129
rect 862 61 872 95
rect 906 61 916 95
rect 862 47 916 61
rect 946 95 1000 177
rect 946 61 956 95
rect 990 61 1000 95
rect 946 47 1000 61
rect 1030 163 1084 177
rect 1030 129 1040 163
rect 1074 129 1084 163
rect 1030 95 1084 129
rect 1030 61 1040 95
rect 1074 61 1084 95
rect 1030 47 1084 61
rect 1114 163 1169 177
rect 1114 129 1124 163
rect 1158 129 1169 163
rect 1114 95 1169 129
rect 1114 61 1124 95
rect 1158 61 1169 95
rect 1114 47 1169 61
<< pdiff >>
rect 27 475 79 494
rect 27 441 35 475
rect 69 441 79 475
rect 27 410 79 441
rect 109 482 161 494
rect 109 448 119 482
rect 153 448 161 482
rect 109 410 161 448
rect 124 381 161 410
rect 336 479 388 497
rect 336 445 344 479
rect 378 445 388 479
rect 124 297 176 381
rect 206 343 258 381
rect 206 309 216 343
rect 250 309 258 343
rect 206 297 258 309
rect 336 297 388 445
rect 418 409 472 497
rect 418 375 428 409
rect 462 375 472 409
rect 418 297 472 375
rect 502 477 556 497
rect 502 443 512 477
rect 546 443 556 477
rect 502 297 556 443
rect 586 341 640 497
rect 586 307 596 341
rect 630 307 640 341
rect 586 297 640 307
rect 670 477 722 497
rect 670 443 680 477
rect 714 443 722 477
rect 670 297 722 443
rect 776 477 832 497
rect 776 443 788 477
rect 822 443 832 477
rect 776 297 832 443
rect 862 409 916 497
rect 862 375 872 409
rect 906 375 916 409
rect 862 341 916 375
rect 862 307 872 341
rect 906 307 916 341
rect 862 297 916 307
rect 946 477 1000 497
rect 946 443 956 477
rect 990 443 1000 477
rect 946 409 1000 443
rect 946 375 956 409
rect 990 375 1000 409
rect 946 341 1000 375
rect 946 307 956 341
rect 990 307 1000 341
rect 946 297 1000 307
rect 1030 477 1084 497
rect 1030 443 1040 477
rect 1074 443 1084 477
rect 1030 409 1084 443
rect 1030 375 1040 409
rect 1074 375 1084 409
rect 1030 297 1084 375
rect 1114 479 1169 497
rect 1114 445 1124 479
rect 1158 445 1169 479
rect 1114 411 1169 445
rect 1114 377 1124 411
rect 1158 377 1169 411
rect 1114 343 1169 377
rect 1114 309 1124 343
rect 1158 309 1169 343
rect 1114 297 1169 309
<< ndiffc >>
rect 43 115 77 149
rect 127 115 161 149
rect 211 115 245 149
rect 328 61 362 95
rect 428 129 462 163
rect 428 61 462 95
rect 512 61 546 95
rect 596 129 630 163
rect 596 61 630 95
rect 680 61 714 95
rect 788 61 822 95
rect 872 129 906 163
rect 872 61 906 95
rect 956 61 990 95
rect 1040 129 1074 163
rect 1040 61 1074 95
rect 1124 129 1158 163
rect 1124 61 1158 95
<< pdiffc >>
rect 35 441 69 475
rect 119 448 153 482
rect 344 445 378 479
rect 216 309 250 343
rect 428 375 462 409
rect 512 443 546 477
rect 596 307 630 341
rect 680 443 714 477
rect 788 443 822 477
rect 872 375 906 409
rect 872 307 906 341
rect 956 443 990 477
rect 956 375 990 409
rect 956 307 990 341
rect 1040 443 1074 477
rect 1040 375 1074 409
rect 1124 445 1158 479
rect 1124 377 1158 411
rect 1124 309 1158 343
<< poly >>
rect 79 494 109 520
rect 388 497 418 523
rect 472 497 502 523
rect 556 497 586 523
rect 640 497 670 523
rect 832 497 862 523
rect 916 497 946 523
rect 1000 497 1030 523
rect 1084 497 1114 523
rect 79 265 109 410
rect 176 381 206 407
rect 176 265 206 297
rect 388 265 418 297
rect 472 265 502 297
rect 556 265 586 297
rect 640 265 670 297
rect 832 265 862 297
rect 916 265 946 297
rect 75 249 129 265
rect 75 215 85 249
rect 119 215 129 249
rect 75 199 129 215
rect 171 249 240 265
rect 171 215 190 249
rect 224 215 240 249
rect 171 199 240 215
rect 350 249 502 265
rect 350 215 360 249
rect 394 215 428 249
rect 462 215 502 249
rect 350 199 502 215
rect 553 249 675 265
rect 553 215 563 249
rect 597 215 631 249
rect 665 215 675 249
rect 553 199 675 215
rect 832 249 946 265
rect 832 215 875 249
rect 909 215 946 249
rect 832 199 946 215
rect 87 177 117 199
rect 171 177 201 199
rect 388 177 418 199
rect 472 177 502 199
rect 556 177 586 199
rect 640 177 670 199
rect 832 177 862 199
rect 916 177 946 199
rect 1000 265 1030 297
rect 1084 265 1114 297
rect 1000 249 1114 265
rect 1000 215 1042 249
rect 1076 215 1114 249
rect 1000 199 1114 215
rect 1000 177 1030 199
rect 1084 177 1114 199
rect 87 67 117 93
rect 171 67 201 93
rect 388 21 418 47
rect 472 21 502 47
rect 556 21 586 47
rect 640 21 670 47
rect 832 21 862 47
rect 916 21 946 47
rect 1000 21 1030 47
rect 1084 21 1114 47
<< polycont >>
rect 85 215 119 249
rect 190 215 224 249
rect 360 215 394 249
rect 428 215 462 249
rect 563 215 597 249
rect 631 215 665 249
rect 875 215 909 249
rect 1042 215 1076 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 482 169 527
rect 103 448 119 482
rect 153 448 169 482
rect 328 479 730 493
rect 328 445 344 479
rect 378 477 730 479
rect 378 459 512 477
rect 378 445 394 459
rect 496 443 512 459
rect 546 443 680 477
rect 714 443 730 477
rect 772 477 998 493
rect 772 443 788 477
rect 822 443 956 477
rect 990 443 998 477
rect 17 411 69 441
rect 17 377 383 411
rect 17 165 51 377
rect 85 249 156 339
rect 199 309 216 343
rect 250 309 315 343
rect 199 305 315 309
rect 119 215 156 249
rect 85 199 156 215
rect 190 249 247 265
rect 224 215 247 249
rect 190 199 247 215
rect 281 249 315 305
rect 349 317 383 377
rect 428 409 462 425
rect 956 409 998 443
rect 462 375 872 409
rect 906 375 922 409
rect 428 359 462 375
rect 864 341 922 375
rect 349 283 546 317
rect 580 307 596 341
rect 630 307 799 341
rect 580 289 799 307
rect 864 307 872 341
rect 906 307 922 341
rect 864 291 922 307
rect 990 375 998 409
rect 956 341 998 375
rect 1032 477 1074 527
rect 1032 443 1040 477
rect 1032 409 1074 443
rect 1032 375 1040 409
rect 1032 359 1074 375
rect 1108 479 1174 493
rect 1108 445 1124 479
rect 1158 445 1174 479
rect 1108 411 1174 445
rect 1108 377 1124 411
rect 1158 377 1174 411
rect 990 325 998 341
rect 1108 343 1174 377
rect 1108 325 1124 343
rect 990 309 1124 325
rect 1158 309 1174 343
rect 990 307 1174 309
rect 956 291 1174 307
rect 512 255 546 283
rect 512 249 681 255
rect 281 215 360 249
rect 394 215 428 249
rect 462 215 478 249
rect 512 215 563 249
rect 597 215 631 249
rect 665 215 681 249
rect 281 165 315 215
rect 715 181 799 289
rect 833 249 992 255
rect 833 215 875 249
rect 909 215 992 249
rect 1026 249 1179 255
rect 1026 215 1042 249
rect 1076 215 1179 249
rect 17 149 93 165
rect 17 115 43 149
rect 77 115 93 149
rect 17 90 93 115
rect 127 149 161 165
rect 127 17 161 115
rect 211 149 315 165
rect 245 131 315 149
rect 412 163 1090 181
rect 245 115 250 131
rect 211 90 250 115
rect 412 129 428 163
rect 462 145 596 163
rect 462 129 478 145
rect 312 95 378 96
rect 312 61 328 95
rect 362 61 378 95
rect 312 17 378 61
rect 412 95 478 129
rect 580 129 596 145
rect 630 145 872 163
rect 630 129 646 145
rect 412 61 428 95
rect 462 61 478 95
rect 412 51 478 61
rect 512 95 546 111
rect 512 17 546 61
rect 580 95 646 129
rect 856 129 872 145
rect 906 145 1040 163
rect 906 129 922 145
rect 580 61 596 95
rect 630 61 646 95
rect 580 51 646 61
rect 680 95 822 111
rect 714 61 788 95
rect 680 17 822 61
rect 856 95 922 129
rect 1024 129 1040 145
rect 1074 129 1090 163
rect 856 61 872 95
rect 906 61 922 95
rect 856 51 922 61
rect 956 95 990 111
rect 956 17 990 61
rect 1024 95 1090 129
rect 1024 61 1040 95
rect 1074 61 1090 95
rect 1024 51 1090 61
rect 1124 163 1179 181
rect 1158 129 1179 163
rect 1124 95 1179 129
rect 1158 61 1179 95
rect 1124 17 1179 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 400 180 0 0 A
port 1 nsew signal input
flabel locali s 673 289 707 323 0 FreeSans 400 180 0 0 Y
port 9 nsew signal output
flabel locali s 857 221 891 255 0 FreeSans 400 180 0 0 B
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4bb_2
rlabel metal1 s 0 -48 1196 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 1196910
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1187586
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.980 0.000 
<< end >>
