magic
tech sky130B
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__via_pol1__example_5595914180854  sky130_fd_pr__via_pol1__example_5595914180854_0
timestamp 1663361622
transform -1 0 16 0 1 31
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180854  sky130_fd_pr__via_pol1__example_5595914180854_1
timestamp 1663361622
transform 1 0 384 0 1 31
box 0 0 1 1
<< properties >>
string GDS_END 35993286
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 35992804
<< end >>
