magic
tech sky130A
magscale 1 2
timestamp 1663361622
use sky130_fd_pr__dfl1__example_55959141808187  sky130_fd_pr__dfl1__example_55959141808187_0
timestamp 1663361622
transform 1 0 -42 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808187  sky130_fd_pr__dfl1__example_55959141808187_1
timestamp 1663361622
transform 1 0 -30 0 1 -2244
box 0 0 1 1
<< properties >>
string GDS_END 258876
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 253940
<< end >>
