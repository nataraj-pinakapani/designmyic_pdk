magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 0 51 169 54 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 51 1 54 4 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel  s 0 46 169 49 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel  s 0 46 1 49 4 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel � s 97 -2 121 24 6 DRN_HVC
port 3 nsew power bidirectional
rlabel 
 s 85 -2 96 9 6 DRN_HVC
port 3 nsew power bidirectional
rlabel 
 s 0 -2 71 14 6 P_CORE
port 4 nsew power bidirectional
rlabel 
 s 97 -2 169 14 6 P_CORE
port 4 nsew power bidirectional
rlabel  s 54 103 115 164 6 P_PAD
port 5 nsew power bidirectional
rlabel � s 47 -2 71 0 8 SRC_BDY_HVC
port 6 nsew ground bidirectional
rlabel 
 s 73 -2 84 1 8 SRC_BDY_HVC
port 6 nsew ground bidirectional
rlabel  s 126 46 169 55 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 126 35 169 38 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 126 50 169 51 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 54 169 55 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 46 169 46 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 126 35 169 38 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 46 47 55 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 35 48 38 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 46 1 46 4 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 50 47 51 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 54 1 55 4 VSSA
port 7 nsew ground bidirectional
rlabel  s 0 35 48 38 6 VSSA
port 7 nsew ground bidirectional
rlabel  s 121 13 169 16 6 VDDA
port 8 nsew power bidirectional
rlabel  s 121 13 169 16 6 VDDA
port 8 nsew power bidirectional
rlabel  s 0 13 48 16 6 VDDA
port 8 nsew power bidirectional
rlabel  s 0 13 48 16 6 VDDA
port 8 nsew power bidirectional
rlabel  s 126 30 169 33 6 VSWITCH
port 9 nsew power bidirectional
rlabel  s 126 30 169 33 6 VSWITCH
port 9 nsew power bidirectional
rlabel  s 0 30 48 33 6 VSWITCH
port 9 nsew power bidirectional
rlabel  s 0 30 48 33 6 VSWITCH
port 9 nsew power bidirectional
rlabel  s 126 62 169 66 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel  s 126 62 169 67 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel  s 0 62 48 66 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel  s 0 62 48 67 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel  s 126 0 169 5 6 VCCHIB
port 11 nsew power bidirectional
rlabel  s 126 0 169 5 6 VCCHIB
port 11 nsew power bidirectional
rlabel  s 0 0 48 5 6 VCCHIB
port 11 nsew power bidirectional
rlabel  s 0 0 48 5 6 VCCHIB
port 11 nsew power bidirectional
rlabel  s 126 68 169 93 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 126 18 169 22 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 121 18 169 22 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 126 68 169 93 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 0 68 48 93 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 0 18 48 22 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 0 18 48 22 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 0 68 48 93 6 VDDIO
port 12 nsew power bidirectional
rlabel  s 126 7 169 11 6 VCCD
port 13 nsew power bidirectional
rlabel  s 126 7 169 12 6 VCCD
port 13 nsew power bidirectional
rlabel  s 0 7 48 11 6 VCCD
port 13 nsew power bidirectional
rlabel  s 0 7 48 12 6 VCCD
port 13 nsew power bidirectional
rlabel  s 128 174 169 198 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 168 190 168 190 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 126 24 169 28 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 126 24 169 28 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 168 174 169 198 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 0 174 48 198 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 1 190 1 190 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 0 24 48 28 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 0 174 1 198 4 VSSIO
port 14 nsew ground bidirectional
rlabel  s 0 24 48 28 6 VSSIO
port 14 nsew ground bidirectional
rlabel  s 126 40 169 44 6 VSSD
port 15 nsew ground bidirectional
rlabel  s 126 40 169 44 6 VSSD
port 15 nsew ground bidirectional
rlabel  s 0 40 48 44 6 VSSD
port 15 nsew ground bidirectional
rlabel  s 0 40 47 44 6 VSSD
port 15 nsew ground bidirectional
rlabel  s 126 56 169 61 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel  s 126 56 169 61 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel  s 0 56 48 61 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel  s 0 56 48 61 6 VSSIO_Q
port 16 nsew ground bidirectional
<< properties >>
string LEFclass PAD POWER
string FIXED_BBOX 0 0 169 198
string LEFview TRUE
<< end >>
