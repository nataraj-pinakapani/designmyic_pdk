magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -66 377 3810 897
<< pwell >>
rect 1022 223 1280 233
rect 1022 217 1848 223
rect 2173 217 3740 283
rect 4 43 3740 217
rect -26 -43 3770 43
<< locali >>
rect 113 333 179 433
rect 389 369 455 471
rect 505 333 578 356
rect 113 299 578 333
rect 505 219 578 299
rect 684 235 750 430
rect 793 235 905 430
rect 2107 235 2327 269
rect 2293 87 2327 235
rect 2809 162 2904 352
rect 2809 87 2843 162
rect 2293 53 2843 87
rect 3652 99 3722 679
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3744 831
rect 124 735 314 741
rect 124 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 314 735
rect 22 541 88 657
rect 124 577 314 701
rect 684 735 863 741
rect 718 701 756 735
rect 790 701 828 735
rect 862 701 863 735
rect 476 611 542 661
rect 476 577 648 611
rect 22 507 578 541
rect 22 263 56 507
rect 527 403 578 507
rect 614 525 648 577
rect 684 561 863 701
rect 899 727 1073 761
rect 899 525 933 727
rect 614 491 933 525
rect 22 219 451 263
rect 22 103 88 219
rect 614 183 648 491
rect 969 381 1003 691
rect 1039 489 1073 727
rect 1109 735 1145 741
rect 1109 701 1110 735
rect 1144 701 1145 735
rect 1109 525 1145 701
rect 1181 727 1419 761
rect 1181 489 1215 727
rect 1039 455 1215 489
rect 1251 419 1306 691
rect 969 347 1167 381
rect 124 113 314 183
rect 124 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 314 113
rect 476 149 648 183
rect 476 99 542 149
rect 684 113 874 199
rect 969 195 1003 347
rect 1101 247 1167 347
rect 1228 285 1306 419
rect 1342 535 1419 727
rect 1699 735 1889 741
rect 1455 671 1661 705
rect 124 73 314 79
rect 684 79 690 113
rect 724 79 762 113
rect 796 79 834 113
rect 868 79 874 113
rect 930 103 1003 195
rect 1040 113 1090 211
rect 684 73 874 79
rect 1040 79 1046 113
rect 1080 79 1090 113
rect 1040 73 1090 79
rect 1126 87 1160 247
rect 1228 211 1262 285
rect 1196 135 1262 211
rect 1342 205 1376 535
rect 1455 355 1489 671
rect 1310 123 1376 205
rect 1412 321 1489 355
rect 1525 535 1591 635
rect 1627 549 1661 671
rect 1699 701 1705 735
rect 1739 701 1777 735
rect 1811 701 1849 735
rect 1883 701 1889 735
rect 1699 585 1889 701
rect 2167 735 2357 751
rect 2167 701 2173 735
rect 2207 701 2245 735
rect 2279 701 2317 735
rect 2351 701 2357 735
rect 2167 657 2357 701
rect 1925 621 2131 655
rect 1925 549 1959 621
rect 2097 587 2436 621
rect 1412 87 1446 321
rect 1525 305 1559 535
rect 1627 515 1959 549
rect 1627 445 1682 515
rect 1995 479 2061 585
rect 1758 445 2061 479
rect 2381 479 2436 587
rect 2472 569 2538 751
rect 2653 735 2843 741
rect 2653 701 2659 735
rect 2693 701 2731 735
rect 2765 701 2803 735
rect 2837 701 2843 735
rect 3163 735 3281 741
rect 3163 701 3169 735
rect 3203 701 3241 735
rect 3275 701 3281 735
rect 2472 535 2584 569
rect 2653 535 2843 701
rect 2879 667 3125 701
rect 2381 445 2514 479
rect 1595 375 2444 409
rect 1595 341 1661 375
rect 1697 305 2305 339
rect 2394 337 2444 375
rect 1525 271 1731 305
rect 1904 291 1970 305
rect 2480 301 2514 445
rect 1525 205 1559 271
rect 1767 255 1833 269
rect 1767 221 1940 255
rect 1482 105 1559 205
rect 1640 113 1830 185
rect 1126 53 1446 87
rect 1640 79 1646 113
rect 1680 79 1718 113
rect 1752 79 1790 113
rect 1824 79 1830 113
rect 1874 103 1940 221
rect 2067 113 2257 199
rect 1640 73 1830 79
rect 2067 79 2073 113
rect 2107 79 2145 113
rect 2179 79 2217 113
rect 2251 79 2257 113
rect 2067 73 2257 79
rect 2419 267 2514 301
rect 2550 422 2584 535
rect 2879 499 2913 667
rect 2742 458 2913 499
rect 2949 435 3015 631
rect 3059 573 3125 667
rect 3163 609 3281 701
rect 3427 735 3616 741
rect 3427 701 3432 735
rect 3466 701 3504 735
rect 3538 701 3576 735
rect 3610 701 3616 735
rect 3059 539 3204 573
rect 2949 422 3117 435
rect 2550 388 3117 422
rect 2419 157 2453 267
rect 2550 231 2584 388
rect 2489 193 2584 231
rect 2620 157 2670 349
rect 2419 123 2670 157
rect 3051 301 3117 388
rect 2940 113 3118 265
rect 3154 165 3204 539
rect 3317 471 3391 629
rect 3427 471 3616 701
rect 3317 335 3383 471
rect 3550 335 3616 435
rect 3317 301 3616 335
rect 3317 165 3383 301
rect 2974 79 3012 113
rect 3046 79 3084 113
rect 2940 73 3118 79
rect 3419 113 3609 265
rect 3419 79 3425 113
rect 3459 79 3497 113
rect 3531 79 3569 113
rect 3603 79 3609 113
rect 3419 73 3609 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3744 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 130 701 164 735
rect 202 701 236 735
rect 274 701 308 735
rect 684 701 718 735
rect 756 701 790 735
rect 828 701 862 735
rect 1110 701 1144 735
rect 130 79 164 113
rect 202 79 236 113
rect 274 79 308 113
rect 690 79 724 113
rect 762 79 796 113
rect 834 79 868 113
rect 1046 79 1080 113
rect 1705 701 1739 735
rect 1777 701 1811 735
rect 1849 701 1883 735
rect 2173 701 2207 735
rect 2245 701 2279 735
rect 2317 701 2351 735
rect 2659 701 2693 735
rect 2731 701 2765 735
rect 2803 701 2837 735
rect 3169 701 3203 735
rect 3241 701 3275 735
rect 1646 79 1680 113
rect 1718 79 1752 113
rect 1790 79 1824 113
rect 2073 79 2107 113
rect 2145 79 2179 113
rect 2217 79 2251 113
rect 3432 701 3466 735
rect 3504 701 3538 735
rect 3576 701 3610 735
rect 2940 79 2974 113
rect 3012 79 3046 113
rect 3084 79 3118 113
rect 3425 79 3459 113
rect 3497 79 3531 113
rect 3569 79 3603 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
<< metal1 >>
rect 0 831 3744 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3744 831
rect 0 791 3744 797
rect 0 735 3744 763
rect 0 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 684 735
rect 718 701 756 735
rect 790 701 828 735
rect 862 701 1110 735
rect 1144 701 1705 735
rect 1739 701 1777 735
rect 1811 701 1849 735
rect 1883 701 2173 735
rect 2207 701 2245 735
rect 2279 701 2317 735
rect 2351 701 2659 735
rect 2693 701 2731 735
rect 2765 701 2803 735
rect 2837 701 3169 735
rect 3203 701 3241 735
rect 3275 701 3432 735
rect 3466 701 3504 735
rect 3538 701 3576 735
rect 3610 701 3744 735
rect 0 689 3744 701
rect 0 113 3744 125
rect 0 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 690 113
rect 724 79 762 113
rect 796 79 834 113
rect 868 79 1046 113
rect 1080 79 1646 113
rect 1680 79 1718 113
rect 1752 79 1790 113
rect 1824 79 2073 113
rect 2107 79 2145 113
rect 2179 79 2217 113
rect 2251 79 2940 113
rect 2974 79 3012 113
rect 3046 79 3084 113
rect 3118 79 3425 113
rect 3459 79 3497 113
rect 3531 79 3569 113
rect 3603 79 3744 113
rect 0 51 3744 79
rect 0 17 3744 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3744 17
rect 0 -23 3744 -17
<< labels >>
rlabel locali s 793 235 905 430 6 CLK
port 1 nsew clock input
rlabel locali s 389 369 455 471 6 D
port 2 nsew signal input
rlabel locali s 684 235 750 430 6 SCD
port 3 nsew signal input
rlabel locali s 505 219 578 299 6 SCE
port 4 nsew signal input
rlabel locali s 113 299 578 333 6 SCE
port 4 nsew signal input
rlabel locali s 505 333 578 356 6 SCE
port 4 nsew signal input
rlabel locali s 113 333 179 433 6 SCE
port 4 nsew signal input
rlabel locali s 2293 53 2843 87 6 SET_B
port 5 nsew signal input
rlabel locali s 2809 87 2843 162 6 SET_B
port 5 nsew signal input
rlabel locali s 2809 162 2904 352 6 SET_B
port 5 nsew signal input
rlabel locali s 2293 87 2327 235 6 SET_B
port 5 nsew signal input
rlabel locali s 2107 235 2327 269 6 SET_B
port 5 nsew signal input
rlabel metal1 s 0 51 3744 125 6 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 -23 3744 23 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s -26 -43 3770 43 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s 4 43 3740 217 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 2173 217 3740 283 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1022 217 1848 223 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1022 223 1280 233 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 791 3744 837 6 VPB
port 8 nsew power bidirectional
rlabel nwell s -66 377 3810 897 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 689 3744 763 6 VPWR
port 9 nsew power bidirectional
rlabel locali s 3652 99 3722 679 6 Q
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3744 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 605350
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hvl/sky130_fd_sc_hvl.gds
string GDS_START 570398
<< end >>
