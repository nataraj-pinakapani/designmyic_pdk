* NGSPICE file created from sky130_fd_pr__rf_npn_11v0_W1p00L1p00.ext - technology: minimum

.subckt sky130_fd_pr__rf_npn_11v0_W1p00L1p00
.ends

