magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect 0 8242 26980 8664
rect 0 302 422 8242
rect 836 1405 26156 7842
rect 26558 302 26980 8242
rect 0 0 26980 302
<< pwell >>
rect 548 7905 26477 8127
rect 548 756 770 7905
rect 26255 756 26477 7905
rect 548 534 26477 756
<< mvpsubdiff >>
rect 574 8033 642 8101
rect 608 7999 642 8033
rect 26176 8067 26211 8101
rect 26245 8067 26280 8101
rect 26314 8067 26349 8101
rect 26383 8067 26451 8101
rect 26176 8033 26451 8067
rect 26176 7999 26211 8033
rect 26245 7999 26280 8033
rect 26314 7999 26349 8033
rect 574 7964 710 7999
rect 608 7930 642 7964
rect 676 7931 710 7964
rect 26108 7965 26349 7999
rect 26108 7931 26143 7965
rect 26177 7931 26212 7965
rect 26246 7931 26281 7965
rect 676 7930 744 7931
rect 574 7896 744 7930
rect 574 7895 710 7896
rect 608 7861 642 7895
rect 676 7862 710 7895
rect 676 7861 744 7862
rect 574 7827 744 7861
rect 574 7826 710 7827
rect 608 7792 642 7826
rect 676 7793 710 7826
rect 676 7792 744 7793
rect 574 7758 744 7792
rect 574 7757 710 7758
rect 608 7723 642 7757
rect 676 7724 710 7757
rect 676 7723 744 7724
rect 574 7689 744 7723
rect 574 7688 710 7689
rect 608 7654 642 7688
rect 676 7655 710 7688
rect 676 7654 744 7655
rect 574 7620 744 7654
rect 574 7619 710 7620
rect 608 7585 642 7619
rect 676 7586 710 7619
rect 676 7585 744 7586
rect 574 7551 744 7585
rect 574 7550 710 7551
rect 608 7516 642 7550
rect 676 7517 710 7550
rect 676 7516 744 7517
rect 574 7482 744 7516
rect 574 7481 710 7482
rect 608 7447 642 7481
rect 676 7448 710 7481
rect 676 7447 744 7448
rect 574 7413 744 7447
rect 574 7412 710 7413
rect 608 7378 642 7412
rect 676 7379 710 7412
rect 676 7378 744 7379
rect 574 7344 744 7378
rect 574 7343 710 7344
rect 608 7309 642 7343
rect 676 7310 710 7343
rect 676 7309 744 7310
rect 574 7275 744 7309
rect 574 7274 710 7275
rect 608 7240 642 7274
rect 676 7241 710 7274
rect 676 7240 744 7241
rect 574 7206 744 7240
rect 574 7205 710 7206
rect 608 7171 642 7205
rect 676 7172 710 7205
rect 676 7171 744 7172
rect 574 7137 744 7171
rect 574 7136 710 7137
rect 608 7102 642 7136
rect 676 7103 710 7136
rect 676 7102 744 7103
rect 574 7068 744 7102
rect 574 7067 710 7068
rect 608 7033 642 7067
rect 676 7034 710 7067
rect 676 7033 744 7034
rect 574 6999 744 7033
rect 574 6998 710 6999
rect 608 6964 642 6998
rect 676 6965 710 6998
rect 676 6964 744 6965
rect 574 6930 744 6964
rect 574 6929 710 6930
rect 608 6895 642 6929
rect 676 6896 710 6929
rect 676 6895 744 6896
rect 574 6861 744 6895
rect 574 6860 710 6861
rect 608 6826 642 6860
rect 676 6827 710 6860
rect 676 6826 744 6827
rect 574 6792 744 6826
rect 574 6791 710 6792
rect 608 6757 642 6791
rect 676 6758 710 6791
rect 676 6757 744 6758
rect 574 6723 744 6757
rect 574 6722 710 6723
rect 608 6688 642 6722
rect 676 6689 710 6722
rect 676 6688 744 6689
rect 574 6654 744 6688
rect 574 6653 710 6654
rect 608 6619 642 6653
rect 676 6620 710 6653
rect 676 6619 744 6620
rect 574 6585 744 6619
rect 574 6584 710 6585
rect 608 6550 642 6584
rect 676 6551 710 6584
rect 676 6550 744 6551
rect 574 6516 744 6550
rect 574 6515 710 6516
rect 608 6481 642 6515
rect 676 6482 710 6515
rect 676 6481 744 6482
rect 574 6447 744 6481
rect 574 6446 710 6447
rect 608 6412 642 6446
rect 676 6413 710 6446
rect 676 6412 744 6413
rect 574 6378 744 6412
rect 574 6377 710 6378
rect 608 6343 642 6377
rect 676 6344 710 6377
rect 676 6343 744 6344
rect 574 6309 744 6343
rect 574 6308 710 6309
rect 608 6274 642 6308
rect 676 6275 710 6308
rect 676 6274 744 6275
rect 574 6240 744 6274
rect 574 6239 710 6240
rect 608 6205 642 6239
rect 676 6206 710 6239
rect 676 6205 744 6206
rect 574 6171 744 6205
rect 574 6170 710 6171
rect 608 6136 642 6170
rect 676 6137 710 6170
rect 676 6136 744 6137
rect 574 6102 744 6136
rect 574 6101 710 6102
rect 608 6067 642 6101
rect 676 6068 710 6101
rect 676 6067 744 6068
rect 574 6033 744 6067
rect 574 6032 710 6033
rect 608 5998 642 6032
rect 676 5999 710 6032
rect 676 5998 744 5999
rect 574 5964 744 5998
rect 574 5963 710 5964
rect 608 5929 642 5963
rect 676 5930 710 5963
rect 676 5929 744 5930
rect 574 5895 744 5929
rect 574 5894 710 5895
rect 608 5860 642 5894
rect 676 5861 710 5894
rect 676 5860 744 5861
rect 574 5826 744 5860
rect 574 5825 710 5826
rect 608 5791 642 5825
rect 676 5792 710 5825
rect 676 5791 744 5792
rect 574 5757 744 5791
rect 574 5756 710 5757
rect 608 5722 642 5756
rect 676 5723 710 5756
rect 676 5722 744 5723
rect 574 5688 744 5722
rect 574 5687 710 5688
rect 608 5653 642 5687
rect 676 5654 710 5687
rect 676 5653 744 5654
rect 574 5619 744 5653
rect 574 5618 710 5619
rect 608 5584 642 5618
rect 676 5585 710 5618
rect 676 5584 744 5585
rect 574 5550 744 5584
rect 574 5549 710 5550
rect 608 5515 642 5549
rect 676 5516 710 5549
rect 676 5515 744 5516
rect 574 5481 744 5515
rect 574 5480 710 5481
rect 608 5446 642 5480
rect 676 5447 710 5480
rect 676 5446 744 5447
rect 574 5412 744 5446
rect 574 5411 710 5412
rect 608 5377 642 5411
rect 676 5378 710 5411
rect 676 5377 744 5378
rect 574 5343 744 5377
rect 574 5342 710 5343
rect 608 5308 642 5342
rect 676 5309 710 5342
rect 676 5308 744 5309
rect 574 5274 744 5308
rect 574 5273 710 5274
rect 676 5240 710 5273
rect 676 5205 744 5240
rect 574 4627 744 4695
rect 608 4593 642 4627
rect 676 4593 710 4627
rect 574 4558 744 4593
rect 608 4524 642 4558
rect 676 4524 710 4558
rect 574 4489 744 4524
rect 608 4455 642 4489
rect 676 4455 710 4489
rect 574 4420 744 4455
rect 608 4386 642 4420
rect 676 4386 710 4420
rect 574 4351 744 4386
rect 608 4317 642 4351
rect 676 4317 710 4351
rect 574 4282 744 4317
rect 608 4248 642 4282
rect 676 4248 710 4282
rect 574 4213 744 4248
rect 608 4179 642 4213
rect 676 4179 710 4213
rect 574 4144 744 4179
rect 608 4110 642 4144
rect 676 4110 710 4144
rect 574 4075 744 4110
rect 608 4041 642 4075
rect 676 4041 710 4075
rect 574 4006 744 4041
rect 608 3972 642 4006
rect 676 3972 710 4006
rect 574 3937 744 3972
rect 608 3903 642 3937
rect 676 3903 710 3937
rect 574 3868 744 3903
rect 608 3834 642 3868
rect 676 3834 710 3868
rect 574 3799 744 3834
rect 608 3765 642 3799
rect 676 3765 710 3799
rect 574 3730 744 3765
rect 608 3696 642 3730
rect 676 3696 710 3730
rect 574 3661 744 3696
rect 608 3627 642 3661
rect 676 3627 710 3661
rect 574 3592 744 3627
rect 608 3558 642 3592
rect 676 3558 710 3592
rect 574 3523 744 3558
rect 608 3489 642 3523
rect 676 3489 710 3523
rect 574 3454 744 3489
rect 608 3420 642 3454
rect 676 3420 710 3454
rect 574 3385 744 3420
rect 608 3351 642 3385
rect 676 3351 710 3385
rect 574 3316 744 3351
rect 608 3282 642 3316
rect 676 3282 710 3316
rect 574 3247 744 3282
rect 608 3213 642 3247
rect 676 3213 710 3247
rect 574 3178 744 3213
rect 26281 2524 26349 2559
rect 26315 2491 26349 2524
rect 26315 2490 26451 2491
rect 26281 2456 26451 2490
rect 26281 2455 26349 2456
rect 26315 2422 26349 2455
rect 26383 2422 26417 2456
rect 26315 2421 26451 2422
rect 26281 2387 26451 2421
rect 26281 2386 26349 2387
rect 26315 2353 26349 2386
rect 26383 2353 26417 2387
rect 26315 2352 26451 2353
rect 26281 2318 26451 2352
rect 26281 2317 26349 2318
rect 26315 2284 26349 2317
rect 26383 2284 26417 2318
rect 26315 2283 26451 2284
rect 26281 2249 26451 2283
rect 26281 2248 26349 2249
rect 26315 2215 26349 2248
rect 26383 2215 26417 2249
rect 26315 2214 26451 2215
rect 26281 2180 26451 2214
rect 26281 2179 26349 2180
rect 26315 2146 26349 2179
rect 26383 2146 26417 2180
rect 26315 2145 26451 2146
rect 26281 2111 26451 2145
rect 26281 2110 26349 2111
rect 26315 2077 26349 2110
rect 26383 2077 26417 2111
rect 26315 2076 26451 2077
rect 26281 2042 26451 2076
rect 26281 2041 26349 2042
rect 26315 2008 26349 2041
rect 26383 2008 26417 2042
rect 26315 2007 26451 2008
rect 26281 1973 26451 2007
rect 26281 1972 26349 1973
rect 26315 1939 26349 1972
rect 26383 1939 26417 1973
rect 26315 1938 26451 1939
rect 26281 1904 26451 1938
rect 26281 1903 26349 1904
rect 26315 1870 26349 1903
rect 26383 1870 26417 1904
rect 26315 1869 26451 1870
rect 26281 1835 26451 1869
rect 26281 1834 26349 1835
rect 26315 1801 26349 1834
rect 26383 1801 26417 1835
rect 26315 1800 26451 1801
rect 26281 1766 26451 1800
rect 26281 1765 26349 1766
rect 26315 1732 26349 1765
rect 26383 1732 26417 1766
rect 26315 1731 26451 1732
rect 26281 1697 26451 1731
rect 26281 1696 26349 1697
rect 26315 1663 26349 1696
rect 26383 1663 26417 1697
rect 26315 1662 26451 1663
rect 26281 1628 26451 1662
rect 26281 1627 26349 1628
rect 26315 1594 26349 1627
rect 26383 1594 26417 1628
rect 26315 1593 26451 1594
rect 26281 1559 26451 1593
rect 26281 1558 26349 1559
rect 26315 1525 26349 1558
rect 26383 1525 26417 1559
rect 26315 1524 26451 1525
rect 26281 1490 26451 1524
rect 26281 1489 26349 1490
rect 26315 1456 26349 1489
rect 26383 1456 26417 1490
rect 26315 1455 26451 1456
rect 26281 1421 26451 1455
rect 26281 1420 26349 1421
rect 26315 1387 26349 1420
rect 26383 1387 26417 1421
rect 26315 1386 26451 1387
rect 26281 1352 26451 1386
rect 26281 1351 26349 1352
rect 26315 1318 26349 1351
rect 26383 1318 26417 1352
rect 26315 1317 26451 1318
rect 26281 1283 26451 1317
rect 26281 1282 26349 1283
rect 26315 1249 26349 1282
rect 26383 1249 26417 1283
rect 26315 1248 26451 1249
rect 26281 1214 26451 1248
rect 26281 1213 26349 1214
rect 26315 1180 26349 1213
rect 26383 1180 26417 1214
rect 26315 1179 26451 1180
rect 26281 1145 26451 1179
rect 26281 1144 26349 1145
rect 26315 1111 26349 1144
rect 26383 1111 26417 1145
rect 26315 1110 26451 1111
rect 26281 1076 26451 1110
rect 26281 1075 26349 1076
rect 26315 1042 26349 1075
rect 26383 1042 26417 1076
rect 26315 1041 26451 1042
rect 26281 1007 26451 1041
rect 26281 1006 26349 1007
rect 26315 973 26349 1006
rect 26383 973 26417 1007
rect 26315 972 26451 973
rect 26281 938 26451 972
rect 26281 937 26349 938
rect 26315 904 26349 937
rect 26383 904 26417 938
rect 26315 903 26451 904
rect 26281 869 26451 903
rect 26281 868 26349 869
rect 26315 835 26349 868
rect 26383 835 26417 869
rect 26315 834 26451 835
rect 26281 800 26451 834
rect 26281 799 26349 800
rect 26315 766 26349 799
rect 26383 766 26417 800
rect 26315 765 26451 766
rect 26281 731 26451 765
rect 26281 730 26349 731
rect 744 696 779 730
rect 813 696 848 730
rect 882 696 917 730
rect 676 662 917 696
rect 26315 697 26349 730
rect 26383 697 26417 731
rect 26315 662 26451 697
rect 676 628 711 662
rect 745 628 780 662
rect 814 628 849 662
rect 574 594 849 628
rect 574 560 642 594
rect 676 560 711 594
rect 745 560 780 594
rect 814 560 849 594
rect 26383 628 26417 662
rect 26383 560 26451 628
<< mvnsubdiff >>
rect 126 8504 249 8538
rect 283 8504 317 8538
rect 126 8470 317 8504
rect 228 8436 317 8470
rect 228 8402 385 8436
rect 296 8368 385 8402
rect 26735 8368 26769 8538
rect 26684 8294 26854 8368
rect 960 7682 1042 7716
rect 1076 7682 1110 7716
rect 960 7648 1110 7682
rect 1062 7614 1110 7648
rect 25964 7615 26032 7716
rect 25964 7614 25998 7615
rect 1062 7580 1178 7614
rect 1130 7546 1178 7580
rect 25896 7581 25998 7614
rect 25896 7547 26032 7581
rect 25896 7546 25930 7547
rect 960 2048 1130 2174
rect 1062 1699 1130 1742
rect 25862 7479 25930 7546
rect 1062 1674 1096 1699
rect 960 1640 1096 1674
rect 994 1631 1096 1640
rect 25814 1665 25862 1699
rect 25814 1631 25930 1665
rect 994 1606 1028 1631
rect 960 1529 1028 1606
rect 25882 1597 25930 1631
rect 25882 1563 26032 1597
rect 25882 1529 25916 1563
rect 25950 1529 26032 1563
rect 364 202 399 236
rect 433 202 468 236
rect 502 202 537 236
rect 571 202 606 236
rect 640 202 675 236
rect 709 202 744 236
rect 778 202 813 236
rect 847 202 882 236
rect 916 202 951 236
rect 985 202 1020 236
rect 1054 202 1089 236
rect 1123 202 1158 236
rect 1192 202 1227 236
rect 1261 202 1296 236
rect 1330 202 1365 236
rect 1399 202 1434 236
rect 1468 202 1503 236
rect 1537 202 1572 236
rect 1606 202 1641 236
rect 1675 202 1710 236
rect 1744 202 1779 236
rect 1813 202 1848 236
rect 1882 202 1917 236
rect 1951 202 1986 236
rect 2020 202 2055 236
rect 2089 202 2124 236
rect 2158 202 2193 236
rect 2227 202 2262 236
rect 2296 202 2331 236
rect 2365 202 2400 236
rect 2434 202 2469 236
rect 2503 202 2538 236
rect 2572 202 2607 236
rect 2641 202 2676 236
rect 2710 202 2745 236
rect 2779 202 2814 236
rect 2848 202 2883 236
rect 2917 202 2952 236
rect 364 168 2952 202
rect 126 134 330 140
rect 364 134 399 168
rect 433 134 468 168
rect 502 134 537 168
rect 571 134 606 168
rect 640 134 675 168
rect 709 134 744 168
rect 778 134 813 168
rect 847 134 882 168
rect 916 134 951 168
rect 985 134 1020 168
rect 1054 134 1089 168
rect 1123 134 1158 168
rect 1192 134 1227 168
rect 1261 134 1296 168
rect 1330 134 1365 168
rect 1399 134 1434 168
rect 1468 134 1503 168
rect 1537 134 1572 168
rect 1606 134 1641 168
rect 1675 134 1710 168
rect 1744 134 1779 168
rect 1813 134 1848 168
rect 1882 134 1917 168
rect 1951 134 1986 168
rect 2020 134 2055 168
rect 2089 134 2124 168
rect 2158 134 2193 168
rect 2227 134 2262 168
rect 2296 134 2331 168
rect 2365 134 2400 168
rect 2434 134 2469 168
rect 2503 134 2538 168
rect 2572 134 2607 168
rect 2641 134 2676 168
rect 2710 134 2745 168
rect 2779 134 2814 168
rect 2848 134 2883 168
rect 2917 134 2952 168
rect 126 100 2952 134
rect 126 66 330 100
rect 364 66 399 100
rect 433 66 468 100
rect 502 66 537 100
rect 571 66 606 100
rect 640 66 675 100
rect 709 66 744 100
rect 778 66 813 100
rect 847 66 882 100
rect 916 66 951 100
rect 985 66 1020 100
rect 1054 66 1089 100
rect 1123 66 1158 100
rect 1192 66 1227 100
rect 1261 66 1296 100
rect 1330 66 1365 100
rect 1399 66 1434 100
rect 1468 66 1503 100
rect 1537 66 1572 100
rect 1606 66 1641 100
rect 1675 66 1710 100
rect 1744 66 1779 100
rect 1813 66 1848 100
rect 1882 66 1917 100
rect 1951 66 1986 100
rect 2020 66 2055 100
rect 2089 66 2124 100
rect 2158 66 2193 100
rect 2227 66 2262 100
rect 2296 66 2331 100
rect 2365 66 2400 100
rect 2434 66 2469 100
rect 2503 66 2538 100
rect 2572 66 2607 100
rect 2641 66 2676 100
rect 2710 66 2745 100
rect 2779 66 2814 100
rect 2848 66 2883 100
rect 2917 66 2952 100
rect 26650 66 26854 100
<< mvpsubdiffcont >>
rect 574 7999 608 8033
rect 642 7999 26176 8101
rect 26211 8067 26245 8101
rect 26280 8067 26314 8101
rect 26349 8067 26383 8101
rect 26211 7999 26245 8033
rect 26280 7999 26314 8033
rect 574 7930 608 7964
rect 642 7930 676 7964
rect 710 7931 26108 7999
rect 26349 7965 26451 8033
rect 26143 7931 26177 7965
rect 26212 7931 26246 7965
rect 574 7861 608 7895
rect 642 7861 676 7895
rect 710 7862 744 7896
rect 574 7792 608 7826
rect 642 7792 676 7826
rect 710 7793 744 7827
rect 574 7723 608 7757
rect 642 7723 676 7757
rect 710 7724 744 7758
rect 574 7654 608 7688
rect 642 7654 676 7688
rect 710 7655 744 7689
rect 574 7585 608 7619
rect 642 7585 676 7619
rect 710 7586 744 7620
rect 574 7516 608 7550
rect 642 7516 676 7550
rect 710 7517 744 7551
rect 574 7447 608 7481
rect 642 7447 676 7481
rect 710 7448 744 7482
rect 574 7378 608 7412
rect 642 7378 676 7412
rect 710 7379 744 7413
rect 574 7309 608 7343
rect 642 7309 676 7343
rect 710 7310 744 7344
rect 574 7240 608 7274
rect 642 7240 676 7274
rect 710 7241 744 7275
rect 574 7171 608 7205
rect 642 7171 676 7205
rect 710 7172 744 7206
rect 574 7102 608 7136
rect 642 7102 676 7136
rect 710 7103 744 7137
rect 574 7033 608 7067
rect 642 7033 676 7067
rect 710 7034 744 7068
rect 574 6964 608 6998
rect 642 6964 676 6998
rect 710 6965 744 6999
rect 574 6895 608 6929
rect 642 6895 676 6929
rect 710 6896 744 6930
rect 574 6826 608 6860
rect 642 6826 676 6860
rect 710 6827 744 6861
rect 574 6757 608 6791
rect 642 6757 676 6791
rect 710 6758 744 6792
rect 574 6688 608 6722
rect 642 6688 676 6722
rect 710 6689 744 6723
rect 574 6619 608 6653
rect 642 6619 676 6653
rect 710 6620 744 6654
rect 574 6550 608 6584
rect 642 6550 676 6584
rect 710 6551 744 6585
rect 574 6481 608 6515
rect 642 6481 676 6515
rect 710 6482 744 6516
rect 574 6412 608 6446
rect 642 6412 676 6446
rect 710 6413 744 6447
rect 574 6343 608 6377
rect 642 6343 676 6377
rect 710 6344 744 6378
rect 574 6274 608 6308
rect 642 6274 676 6308
rect 710 6275 744 6309
rect 574 6205 608 6239
rect 642 6205 676 6239
rect 710 6206 744 6240
rect 574 6136 608 6170
rect 642 6136 676 6170
rect 710 6137 744 6171
rect 574 6067 608 6101
rect 642 6067 676 6101
rect 710 6068 744 6102
rect 574 5998 608 6032
rect 642 5998 676 6032
rect 710 5999 744 6033
rect 574 5929 608 5963
rect 642 5929 676 5963
rect 710 5930 744 5964
rect 574 5860 608 5894
rect 642 5860 676 5894
rect 710 5861 744 5895
rect 574 5791 608 5825
rect 642 5791 676 5825
rect 710 5792 744 5826
rect 574 5722 608 5756
rect 642 5722 676 5756
rect 710 5723 744 5757
rect 574 5653 608 5687
rect 642 5653 676 5687
rect 710 5654 744 5688
rect 574 5584 608 5618
rect 642 5584 676 5618
rect 710 5585 744 5619
rect 574 5515 608 5549
rect 642 5515 676 5549
rect 710 5516 744 5550
rect 574 5446 608 5480
rect 642 5446 676 5480
rect 710 5447 744 5481
rect 574 5377 608 5411
rect 642 5377 676 5411
rect 710 5378 744 5412
rect 574 5308 608 5342
rect 642 5308 676 5342
rect 710 5309 744 5343
rect 574 5205 676 5273
rect 710 5240 744 5274
rect 574 4695 744 5205
rect 574 4593 608 4627
rect 642 4593 676 4627
rect 710 4593 744 4627
rect 574 4524 608 4558
rect 642 4524 676 4558
rect 710 4524 744 4558
rect 574 4455 608 4489
rect 642 4455 676 4489
rect 710 4455 744 4489
rect 574 4386 608 4420
rect 642 4386 676 4420
rect 710 4386 744 4420
rect 574 4317 608 4351
rect 642 4317 676 4351
rect 710 4317 744 4351
rect 574 4248 608 4282
rect 642 4248 676 4282
rect 710 4248 744 4282
rect 574 4179 608 4213
rect 642 4179 676 4213
rect 710 4179 744 4213
rect 574 4110 608 4144
rect 642 4110 676 4144
rect 710 4110 744 4144
rect 574 4041 608 4075
rect 642 4041 676 4075
rect 710 4041 744 4075
rect 574 3972 608 4006
rect 642 3972 676 4006
rect 710 3972 744 4006
rect 574 3903 608 3937
rect 642 3903 676 3937
rect 710 3903 744 3937
rect 574 3834 608 3868
rect 642 3834 676 3868
rect 710 3834 744 3868
rect 574 3765 608 3799
rect 642 3765 676 3799
rect 710 3765 744 3799
rect 574 3696 608 3730
rect 642 3696 676 3730
rect 710 3696 744 3730
rect 574 3627 608 3661
rect 642 3627 676 3661
rect 710 3627 744 3661
rect 574 3558 608 3592
rect 642 3558 676 3592
rect 710 3558 744 3592
rect 574 3489 608 3523
rect 642 3489 676 3523
rect 710 3489 744 3523
rect 574 3420 608 3454
rect 642 3420 676 3454
rect 710 3420 744 3454
rect 574 3351 608 3385
rect 642 3351 676 3385
rect 710 3351 744 3385
rect 574 3282 608 3316
rect 642 3282 676 3316
rect 710 3282 744 3316
rect 574 3213 608 3247
rect 642 3213 676 3247
rect 710 3213 744 3247
rect 574 696 744 3178
rect 26281 2559 26451 7965
rect 26281 2490 26315 2524
rect 26349 2491 26451 2559
rect 26281 2421 26315 2455
rect 26349 2422 26383 2456
rect 26417 2422 26451 2456
rect 26281 2352 26315 2386
rect 26349 2353 26383 2387
rect 26417 2353 26451 2387
rect 26281 2283 26315 2317
rect 26349 2284 26383 2318
rect 26417 2284 26451 2318
rect 26281 2214 26315 2248
rect 26349 2215 26383 2249
rect 26417 2215 26451 2249
rect 26281 2145 26315 2179
rect 26349 2146 26383 2180
rect 26417 2146 26451 2180
rect 26281 2076 26315 2110
rect 26349 2077 26383 2111
rect 26417 2077 26451 2111
rect 26281 2007 26315 2041
rect 26349 2008 26383 2042
rect 26417 2008 26451 2042
rect 26281 1938 26315 1972
rect 26349 1939 26383 1973
rect 26417 1939 26451 1973
rect 26281 1869 26315 1903
rect 26349 1870 26383 1904
rect 26417 1870 26451 1904
rect 26281 1800 26315 1834
rect 26349 1801 26383 1835
rect 26417 1801 26451 1835
rect 26281 1731 26315 1765
rect 26349 1732 26383 1766
rect 26417 1732 26451 1766
rect 26281 1662 26315 1696
rect 26349 1663 26383 1697
rect 26417 1663 26451 1697
rect 26281 1593 26315 1627
rect 26349 1594 26383 1628
rect 26417 1594 26451 1628
rect 26281 1524 26315 1558
rect 26349 1525 26383 1559
rect 26417 1525 26451 1559
rect 26281 1455 26315 1489
rect 26349 1456 26383 1490
rect 26417 1456 26451 1490
rect 26281 1386 26315 1420
rect 26349 1387 26383 1421
rect 26417 1387 26451 1421
rect 26281 1317 26315 1351
rect 26349 1318 26383 1352
rect 26417 1318 26451 1352
rect 26281 1248 26315 1282
rect 26349 1249 26383 1283
rect 26417 1249 26451 1283
rect 26281 1179 26315 1213
rect 26349 1180 26383 1214
rect 26417 1180 26451 1214
rect 26281 1110 26315 1144
rect 26349 1111 26383 1145
rect 26417 1111 26451 1145
rect 26281 1041 26315 1075
rect 26349 1042 26383 1076
rect 26417 1042 26451 1076
rect 26281 972 26315 1006
rect 26349 973 26383 1007
rect 26417 973 26451 1007
rect 26281 903 26315 937
rect 26349 904 26383 938
rect 26417 904 26451 938
rect 26281 834 26315 868
rect 26349 835 26383 869
rect 26417 835 26451 869
rect 26281 765 26315 799
rect 26349 766 26383 800
rect 26417 766 26451 800
rect 779 696 813 730
rect 848 696 882 730
rect 574 628 676 696
rect 917 662 26315 730
rect 26349 697 26383 731
rect 26417 697 26451 731
rect 711 628 745 662
rect 780 628 814 662
rect 642 560 676 594
rect 711 560 745 594
rect 780 560 814 594
rect 849 560 26383 662
rect 26417 628 26451 662
<< mvnsubdiffcont >>
rect 249 8504 283 8538
rect 126 8402 228 8470
rect 317 8436 26735 8538
rect 126 236 296 8402
rect 385 8368 26735 8436
rect 1042 7682 1076 7716
rect 960 7580 1062 7648
rect 1110 7614 25964 7716
rect 960 2174 1130 7580
rect 1178 7546 25896 7614
rect 25998 7581 26032 7615
rect 960 1742 1130 2048
rect 960 1674 1062 1742
rect 25930 7479 26032 7547
rect 960 1606 994 1640
rect 1096 1631 25814 1699
rect 25862 1665 26032 7479
rect 1028 1529 25882 1631
rect 25930 1597 26032 1665
rect 25916 1529 25950 1563
rect 26684 236 26854 8294
rect 126 140 364 236
rect 399 202 433 236
rect 468 202 502 236
rect 537 202 571 236
rect 606 202 640 236
rect 675 202 709 236
rect 744 202 778 236
rect 813 202 847 236
rect 882 202 916 236
rect 951 202 985 236
rect 1020 202 1054 236
rect 1089 202 1123 236
rect 1158 202 1192 236
rect 1227 202 1261 236
rect 1296 202 1330 236
rect 1365 202 1399 236
rect 1434 202 1468 236
rect 1503 202 1537 236
rect 1572 202 1606 236
rect 1641 202 1675 236
rect 1710 202 1744 236
rect 1779 202 1813 236
rect 1848 202 1882 236
rect 1917 202 1951 236
rect 1986 202 2020 236
rect 2055 202 2089 236
rect 2124 202 2158 236
rect 2193 202 2227 236
rect 2262 202 2296 236
rect 2331 202 2365 236
rect 2400 202 2434 236
rect 2469 202 2503 236
rect 2538 202 2572 236
rect 2607 202 2641 236
rect 2676 202 2710 236
rect 2745 202 2779 236
rect 2814 202 2848 236
rect 2883 202 2917 236
rect 330 134 364 140
rect 399 134 433 168
rect 468 134 502 168
rect 537 134 571 168
rect 606 134 640 168
rect 675 134 709 168
rect 744 134 778 168
rect 813 134 847 168
rect 882 134 916 168
rect 951 134 985 168
rect 1020 134 1054 168
rect 1089 134 1123 168
rect 1158 134 1192 168
rect 1227 134 1261 168
rect 1296 134 1330 168
rect 1365 134 1399 168
rect 1434 134 1468 168
rect 1503 134 1537 168
rect 1572 134 1606 168
rect 1641 134 1675 168
rect 1710 134 1744 168
rect 1779 134 1813 168
rect 1848 134 1882 168
rect 1917 134 1951 168
rect 1986 134 2020 168
rect 2055 134 2089 168
rect 2124 134 2158 168
rect 2193 134 2227 168
rect 2262 134 2296 168
rect 2331 134 2365 168
rect 2400 134 2434 168
rect 2469 134 2503 168
rect 2538 134 2572 168
rect 2607 134 2641 168
rect 2676 134 2710 168
rect 2745 134 2779 168
rect 2814 134 2848 168
rect 2883 134 2917 168
rect 2952 100 26854 236
rect 330 66 364 100
rect 399 66 433 100
rect 468 66 502 100
rect 537 66 571 100
rect 606 66 640 100
rect 675 66 709 100
rect 744 66 778 100
rect 813 66 847 100
rect 882 66 916 100
rect 951 66 985 100
rect 1020 66 1054 100
rect 1089 66 1123 100
rect 1158 66 1192 100
rect 1227 66 1261 100
rect 1296 66 1330 100
rect 1365 66 1399 100
rect 1434 66 1468 100
rect 1503 66 1537 100
rect 1572 66 1606 100
rect 1641 66 1675 100
rect 1710 66 1744 100
rect 1779 66 1813 100
rect 1848 66 1882 100
rect 1917 66 1951 100
rect 1986 66 2020 100
rect 2055 66 2089 100
rect 2124 66 2158 100
rect 2193 66 2227 100
rect 2262 66 2296 100
rect 2331 66 2365 100
rect 2400 66 2434 100
rect 2469 66 2503 100
rect 2538 66 2572 100
rect 2607 66 2641 100
rect 2676 66 2710 100
rect 2745 66 2779 100
rect 2814 66 2848 100
rect 2883 66 2917 100
rect 2952 66 26650 100
<< locali >>
rect 126 8504 249 8538
rect 283 8504 317 8538
rect 126 8490 317 8504
rect 116 8484 317 8490
rect 26735 8490 26769 8538
rect 116 8470 194 8484
rect 116 8412 126 8470
rect 228 8450 267 8484
rect 301 8450 317 8484
rect 228 8436 317 8450
rect 228 8412 385 8436
rect 116 1250 122 8412
rect 228 8402 267 8412
rect 301 8378 340 8412
rect 374 8378 385 8412
rect 26735 8452 26864 8490
rect 26735 8418 26752 8452
rect 26786 8418 26824 8452
rect 26858 8418 26864 8452
rect 296 8368 385 8378
rect 26735 8372 26864 8418
rect 26735 8368 26752 8372
rect 296 8340 4354 8368
rect 300 8306 339 8340
rect 373 8306 412 8340
rect 446 8306 485 8340
rect 519 8306 558 8340
rect 592 8306 631 8340
rect 665 8306 704 8340
rect 738 8306 777 8340
rect 811 8306 850 8340
rect 884 8306 923 8340
rect 957 8306 996 8340
rect 1030 8306 1069 8340
rect 1103 8306 1142 8340
rect 1176 8306 1215 8340
rect 1249 8306 1288 8340
rect 1322 8306 1361 8340
rect 1395 8306 1434 8340
rect 1468 8306 1507 8340
rect 1541 8306 1580 8340
rect 1614 8306 1653 8340
rect 1687 8306 1726 8340
rect 1760 8306 1799 8340
rect 1833 8306 1872 8340
rect 1906 8306 1945 8340
rect 1979 8306 2018 8340
rect 2052 8306 2091 8340
rect 2125 8306 2164 8340
rect 2198 8306 2237 8340
rect 2271 8306 2310 8340
rect 2344 8306 2383 8340
rect 2417 8306 2456 8340
rect 2490 8306 2529 8340
rect 2563 8306 2602 8340
rect 2636 8306 2675 8340
rect 2709 8306 2748 8340
rect 2782 8306 2821 8340
rect 2855 8306 2894 8340
rect 2928 8306 2967 8340
rect 3001 8306 3040 8340
rect 3074 8306 3113 8340
rect 3147 8306 3186 8340
rect 3220 8306 3259 8340
rect 3293 8306 3332 8340
rect 3366 8306 3405 8340
rect 3439 8306 3478 8340
rect 3512 8306 3551 8340
rect 3585 8306 3624 8340
rect 3658 8306 3697 8340
rect 3731 8306 3770 8340
rect 3804 8306 3843 8340
rect 3877 8306 3916 8340
rect 3950 8306 3989 8340
rect 4023 8306 4062 8340
rect 4096 8306 4135 8340
rect 4169 8306 4208 8340
rect 4242 8306 4281 8340
rect 4315 8306 4354 8340
rect 26636 8338 26680 8368
rect 26714 8338 26752 8368
rect 26786 8338 26824 8372
rect 26858 8338 26864 8372
rect 26636 8306 26864 8338
rect 300 8300 26864 8306
rect 300 1322 306 8300
rect 26674 8294 26864 8300
rect 26674 8292 26684 8294
rect 26854 8292 26864 8294
rect 26674 8258 26680 8292
rect 26858 8258 26864 8292
rect 26674 8212 26684 8258
rect 26854 8212 26864 8258
rect 26674 8178 26680 8212
rect 26858 8178 26864 8212
rect 26674 8133 26684 8178
rect 26854 8133 26864 8178
rect 296 1283 306 1322
rect 116 1211 126 1250
rect 300 1249 306 1283
rect 116 1177 122 1211
rect 296 1210 306 1249
rect 116 1138 126 1177
rect 300 1176 306 1210
rect 116 1104 122 1138
rect 296 1137 306 1176
rect 116 1065 126 1104
rect 300 1103 306 1137
rect 116 1031 122 1065
rect 296 1064 306 1103
rect 116 992 126 1031
rect 300 1030 306 1064
rect 116 958 122 992
rect 296 991 306 1030
rect 116 919 126 958
rect 300 957 306 991
rect 116 885 122 919
rect 296 918 306 957
rect 116 846 126 885
rect 300 884 306 918
rect 116 812 122 846
rect 296 845 306 884
rect 116 773 126 812
rect 300 811 306 845
rect 116 739 122 773
rect 296 772 306 811
rect 116 700 126 739
rect 300 738 306 772
rect 116 666 122 700
rect 296 699 306 738
rect 116 627 126 666
rect 300 665 306 699
rect 116 593 122 627
rect 296 626 306 665
rect 116 554 126 593
rect 300 592 306 626
rect 116 520 122 554
rect 296 553 306 592
rect 116 481 126 520
rect 300 519 306 553
rect 564 8105 26461 8111
rect 564 8033 642 8105
rect 676 8101 715 8105
rect 749 8101 788 8105
rect 822 8101 861 8105
rect 564 4615 570 8033
rect 26383 8033 26461 8105
rect 26455 7999 26461 8033
rect 676 7961 710 7999
rect 26311 7965 26349 7999
rect 748 7927 787 7931
rect 821 7927 860 7931
rect 894 7927 933 7931
rect 26451 7959 26461 7999
rect 748 7921 26281 7927
rect 26455 7925 26461 7959
rect 748 4687 754 7921
rect 26271 7887 26281 7921
rect 26271 7853 26277 7887
rect 26451 7885 26461 7925
rect 26271 7813 26281 7853
rect 26455 7851 26461 7885
rect 26271 7779 26277 7813
rect 26451 7811 26461 7851
rect 26271 7739 26281 7779
rect 26455 7777 26461 7811
rect 676 4648 754 4687
rect 676 4627 714 4648
rect 564 4593 574 4615
rect 608 4593 642 4615
rect 676 4593 710 4627
rect 748 4614 754 4648
rect 744 4593 754 4614
rect 564 4576 754 4593
rect 564 4542 570 4576
rect 604 4558 642 4576
rect 676 4575 754 4576
rect 676 4558 714 4575
rect 564 4524 574 4542
rect 608 4524 642 4558
rect 676 4524 710 4558
rect 748 4541 754 4575
rect 744 4524 754 4541
rect 564 4503 754 4524
rect 564 4469 570 4503
rect 604 4489 642 4503
rect 676 4502 754 4503
rect 676 4489 714 4502
rect 564 4455 574 4469
rect 608 4455 642 4489
rect 676 4455 710 4489
rect 748 4468 754 4502
rect 744 4455 754 4468
rect 564 4430 754 4455
rect 564 4396 570 4430
rect 604 4420 642 4430
rect 676 4429 754 4430
rect 676 4420 714 4429
rect 564 4386 574 4396
rect 608 4386 642 4420
rect 676 4386 710 4420
rect 748 4395 754 4429
rect 744 4386 754 4395
rect 564 4357 754 4386
rect 564 4323 570 4357
rect 604 4351 642 4357
rect 676 4356 754 4357
rect 676 4351 714 4356
rect 564 4317 574 4323
rect 608 4317 642 4351
rect 676 4317 710 4351
rect 748 4322 754 4356
rect 744 4317 754 4322
rect 564 4284 754 4317
rect 564 4250 570 4284
rect 604 4282 642 4284
rect 676 4283 754 4284
rect 676 4282 714 4283
rect 564 4248 574 4250
rect 608 4248 642 4282
rect 676 4248 710 4282
rect 748 4249 754 4283
rect 744 4248 754 4249
rect 564 4213 754 4248
rect 564 4211 574 4213
rect 564 4177 570 4211
rect 608 4179 642 4213
rect 676 4179 710 4213
rect 744 4210 754 4213
rect 604 4177 642 4179
rect 676 4177 714 4179
rect 564 4176 714 4177
rect 748 4176 754 4210
rect 564 4144 754 4176
rect 564 4138 574 4144
rect 564 4104 570 4138
rect 608 4110 642 4144
rect 676 4110 710 4144
rect 744 4137 754 4144
rect 604 4104 642 4110
rect 676 4104 714 4110
rect 564 4103 714 4104
rect 748 4103 754 4137
rect 564 4075 754 4103
rect 564 4065 574 4075
rect 564 4031 570 4065
rect 608 4041 642 4075
rect 676 4041 710 4075
rect 744 4064 754 4075
rect 604 4031 642 4041
rect 676 4031 714 4041
rect 564 4030 714 4031
rect 748 4030 754 4064
rect 564 4006 754 4030
rect 564 3992 574 4006
rect 564 3958 570 3992
rect 608 3972 642 4006
rect 676 3972 710 4006
rect 744 3991 754 4006
rect 604 3958 642 3972
rect 676 3958 714 3972
rect 564 3957 714 3958
rect 748 3957 754 3991
rect 564 3937 754 3957
rect 564 3919 574 3937
rect 564 3885 570 3919
rect 608 3903 642 3937
rect 676 3903 710 3937
rect 744 3918 754 3937
rect 604 3885 642 3903
rect 676 3885 714 3903
rect 564 3884 714 3885
rect 748 3884 754 3918
rect 564 3868 754 3884
rect 564 3846 574 3868
rect 564 3812 570 3846
rect 608 3834 642 3868
rect 676 3834 710 3868
rect 744 3845 754 3868
rect 604 3812 642 3834
rect 676 3812 714 3834
rect 564 3811 714 3812
rect 748 3811 754 3845
rect 564 3799 754 3811
rect 564 3773 574 3799
rect 564 3739 570 3773
rect 608 3765 642 3799
rect 676 3765 710 3799
rect 744 3772 754 3799
rect 604 3739 642 3765
rect 676 3739 714 3765
rect 564 3738 714 3739
rect 748 3738 754 3772
rect 564 3730 754 3738
rect 564 3700 574 3730
rect 564 3666 570 3700
rect 608 3696 642 3730
rect 676 3696 710 3730
rect 744 3699 754 3730
rect 604 3666 642 3696
rect 676 3666 714 3696
rect 564 3665 714 3666
rect 748 3665 754 3699
rect 564 3661 754 3665
rect 564 3627 574 3661
rect 608 3627 642 3661
rect 676 3627 710 3661
rect 744 3627 754 3661
rect 564 3593 570 3627
rect 604 3593 642 3627
rect 676 3626 754 3627
rect 676 3593 714 3626
rect 564 3592 714 3593
rect 748 3592 754 3626
rect 564 3558 574 3592
rect 608 3558 642 3592
rect 676 3558 710 3592
rect 744 3558 754 3592
rect 564 3554 754 3558
rect 564 3520 570 3554
rect 604 3523 642 3554
rect 676 3553 754 3554
rect 676 3523 714 3553
rect 564 3489 574 3520
rect 608 3489 642 3523
rect 676 3489 710 3523
rect 748 3519 754 3553
rect 744 3489 754 3519
rect 564 3481 754 3489
rect 564 3447 570 3481
rect 604 3454 642 3481
rect 676 3480 754 3481
rect 676 3454 714 3480
rect 564 3420 574 3447
rect 608 3420 642 3454
rect 676 3420 710 3454
rect 748 3446 754 3480
rect 744 3420 754 3446
rect 564 3408 754 3420
rect 564 3374 570 3408
rect 604 3385 642 3408
rect 676 3407 754 3408
rect 676 3385 714 3407
rect 564 3351 574 3374
rect 608 3351 642 3385
rect 676 3351 710 3385
rect 748 3373 754 3407
rect 744 3351 754 3373
rect 564 3335 754 3351
rect 564 3301 570 3335
rect 604 3316 642 3335
rect 676 3334 754 3335
rect 676 3316 714 3334
rect 564 3282 574 3301
rect 608 3282 642 3316
rect 676 3282 710 3316
rect 748 3300 754 3334
rect 744 3282 754 3300
rect 564 3262 754 3282
rect 564 3228 570 3262
rect 604 3247 642 3262
rect 676 3261 754 3262
rect 676 3247 714 3261
rect 564 3213 574 3228
rect 608 3213 642 3247
rect 676 3213 710 3247
rect 748 3227 754 3261
rect 744 3213 754 3227
rect 564 3189 754 3213
rect 564 3155 570 3189
rect 604 3178 642 3189
rect 676 3188 754 3189
rect 676 3178 714 3188
rect 564 3116 574 3155
rect 748 3154 754 3188
rect 564 3082 570 3116
rect 744 3115 754 3154
rect 564 3043 574 3082
rect 748 3081 754 3115
rect 564 3009 570 3043
rect 744 3042 754 3081
rect 564 2970 574 3009
rect 748 3008 754 3042
rect 564 2936 570 2970
rect 744 2969 754 3008
rect 564 2897 574 2936
rect 748 2935 754 2969
rect 564 2863 570 2897
rect 744 2896 754 2935
rect 564 2824 574 2863
rect 748 2862 754 2896
rect 564 2790 570 2824
rect 744 2823 754 2862
rect 564 2751 574 2790
rect 748 2789 754 2823
rect 564 2717 570 2751
rect 744 2750 754 2789
rect 564 2678 574 2717
rect 748 2716 754 2750
rect 564 2644 570 2678
rect 744 2677 754 2716
rect 564 2605 574 2644
rect 748 2643 754 2677
rect 564 2571 570 2605
rect 744 2604 754 2643
rect 564 2532 574 2571
rect 748 2570 754 2604
rect 564 2498 570 2532
rect 744 2531 754 2570
rect 564 2459 574 2498
rect 748 2497 754 2531
rect 564 2425 570 2459
rect 744 2458 754 2497
rect 564 2386 574 2425
rect 748 2424 754 2458
rect 564 2352 570 2386
rect 744 2385 754 2424
rect 564 2313 574 2352
rect 748 2351 754 2385
rect 564 2279 570 2313
rect 744 2312 754 2351
rect 564 2240 574 2279
rect 748 2278 754 2312
rect 564 2206 570 2240
rect 744 2239 754 2278
rect 564 2167 574 2206
rect 748 2205 754 2239
rect 564 2133 570 2167
rect 744 2166 754 2205
rect 564 2094 574 2133
rect 748 2132 754 2166
rect 564 2060 570 2094
rect 744 2093 754 2132
rect 564 2021 574 2060
rect 748 2059 754 2093
rect 564 1987 570 2021
rect 744 2020 754 2059
rect 564 1948 574 1987
rect 748 1986 754 2020
rect 564 1914 570 1948
rect 744 1947 754 1986
rect 564 1875 574 1914
rect 748 1913 754 1947
rect 564 1841 570 1875
rect 744 1874 754 1913
rect 564 1802 574 1841
rect 748 1840 754 1874
rect 564 1768 570 1802
rect 744 1801 754 1840
rect 564 1729 574 1768
rect 748 1767 754 1801
rect 564 1695 570 1729
rect 744 1728 754 1767
rect 564 1656 574 1695
rect 748 1694 754 1728
rect 564 1622 570 1656
rect 744 1655 754 1694
rect 564 1583 574 1622
rect 748 1621 754 1655
rect 564 1549 570 1583
rect 744 1582 754 1621
rect 564 1510 574 1549
rect 748 1548 754 1582
rect 564 1476 570 1510
rect 744 1509 754 1548
rect 950 7719 26063 7725
rect 950 7685 1028 7719
rect 1062 7716 1101 7719
rect 1135 7716 1174 7719
rect 1208 7716 1247 7719
rect 1281 7716 1320 7719
rect 1354 7716 1393 7719
rect 1427 7716 1466 7719
rect 1500 7716 1539 7719
rect 1573 7716 1612 7719
rect 1646 7716 1685 7719
rect 1719 7716 1758 7719
rect 1792 7716 1831 7719
rect 1076 7685 1101 7716
rect 950 7682 1042 7685
rect 1076 7682 1110 7685
rect 950 7648 1110 7682
rect 950 7647 960 7648
rect 1062 7647 1110 7648
rect 950 4517 956 7647
rect 1062 7613 1101 7647
rect 1135 7613 1174 7614
rect 25985 7647 26063 7719
rect 25985 7615 26023 7647
rect 25985 7613 25998 7615
rect 26057 7613 26063 7647
rect 1062 7580 1178 7613
rect 1130 7575 1178 7580
rect 1134 7541 1173 7575
rect 25913 7581 25998 7613
rect 26032 7581 26063 7613
rect 25913 7573 26063 7581
rect 25913 7547 25951 7573
rect 25985 7547 26023 7573
rect 1207 7541 1246 7546
rect 1280 7541 1319 7546
rect 1353 7541 1392 7546
rect 1426 7541 1465 7546
rect 1499 7541 1538 7546
rect 1572 7541 1611 7546
rect 1645 7541 1684 7546
rect 1718 7541 1757 7546
rect 1791 7541 1830 7546
rect 1864 7541 1903 7546
rect 25913 7541 25930 7547
rect 1134 7535 25930 7541
rect 26057 7539 26063 7573
rect 1134 4589 1140 7535
rect 1130 4550 1140 4589
rect 950 4478 960 4517
rect 1134 4516 1140 4550
rect 950 4444 956 4478
rect 1130 4477 1140 4516
rect 950 4405 960 4444
rect 1134 4443 1140 4477
rect 950 4371 956 4405
rect 1130 4404 1140 4443
rect 950 4332 960 4371
rect 1134 4370 1140 4404
rect 950 4298 956 4332
rect 1130 4331 1140 4370
rect 950 4259 960 4298
rect 1134 4297 1140 4331
rect 950 4225 956 4259
rect 1130 4258 1140 4297
rect 950 4186 960 4225
rect 1134 4224 1140 4258
rect 950 4152 956 4186
rect 1130 4185 1140 4224
rect 950 4113 960 4152
rect 1134 4151 1140 4185
rect 950 4079 956 4113
rect 1130 4112 1140 4151
rect 950 4040 960 4079
rect 1134 4078 1140 4112
rect 950 4006 956 4040
rect 1130 4039 1140 4078
rect 950 3967 960 4006
rect 1134 4005 1140 4039
rect 950 3933 956 3967
rect 1130 3966 1140 4005
rect 950 3894 960 3933
rect 1134 3932 1140 3966
rect 950 3860 956 3894
rect 1130 3893 1140 3932
rect 950 3821 960 3860
rect 1134 3859 1140 3893
rect 950 3787 956 3821
rect 1130 3820 1140 3859
rect 950 3748 960 3787
rect 1134 3786 1140 3820
rect 950 3714 956 3748
rect 1130 3747 1140 3786
rect 950 3675 960 3714
rect 1134 3713 1140 3747
rect 950 3641 956 3675
rect 1130 3674 1140 3713
rect 950 3602 960 3641
rect 1134 3640 1140 3674
rect 950 3568 956 3602
rect 1130 3601 1140 3640
rect 950 3529 960 3568
rect 1134 3567 1140 3601
rect 950 3495 956 3529
rect 1130 3528 1140 3567
rect 950 3456 960 3495
rect 1134 3494 1140 3528
rect 950 3422 956 3456
rect 1130 3455 1140 3494
rect 950 3383 960 3422
rect 1134 3421 1140 3455
rect 950 3349 956 3383
rect 1130 3382 1140 3421
rect 950 3310 960 3349
rect 1134 3348 1140 3382
rect 950 3276 956 3310
rect 1130 3309 1140 3348
rect 950 3237 960 3276
rect 1134 3275 1140 3309
rect 950 3203 956 3237
rect 1130 3236 1140 3275
rect 950 3164 960 3203
rect 1134 3202 1140 3236
rect 950 3130 956 3164
rect 1130 3163 1140 3202
rect 950 3091 960 3130
rect 1134 3129 1140 3163
rect 950 3057 956 3091
rect 1130 3090 1140 3129
rect 950 3018 960 3057
rect 1134 3056 1140 3090
rect 950 2984 956 3018
rect 1130 3017 1140 3056
rect 950 2945 960 2984
rect 1134 2983 1140 3017
rect 950 2911 956 2945
rect 1130 2944 1140 2983
rect 950 2872 960 2911
rect 1134 2910 1140 2944
rect 950 2838 956 2872
rect 1130 2871 1140 2910
rect 950 2799 960 2838
rect 1134 2837 1140 2871
rect 950 2765 956 2799
rect 1130 2798 1140 2837
rect 950 2726 960 2765
rect 1134 2764 1140 2798
rect 950 2692 956 2726
rect 1130 2725 1140 2764
rect 950 2653 960 2692
rect 1134 2691 1140 2725
rect 950 2619 956 2653
rect 1130 2652 1140 2691
rect 950 2580 960 2619
rect 1134 2618 1140 2652
rect 950 2546 956 2580
rect 1130 2579 1140 2618
rect 950 2507 960 2546
rect 1134 2545 1140 2579
rect 950 2473 956 2507
rect 1130 2506 1140 2545
rect 950 2434 960 2473
rect 1134 2472 1140 2506
rect 950 2400 956 2434
rect 1130 2433 1140 2472
rect 950 2361 960 2400
rect 1134 2399 1140 2433
rect 950 2327 956 2361
rect 1130 2360 1140 2399
rect 950 2288 960 2327
rect 1134 2326 1140 2360
rect 950 2254 956 2288
rect 1130 2287 1140 2326
rect 950 2215 960 2254
rect 1134 2253 1140 2287
rect 950 2181 956 2215
rect 1130 2214 1140 2253
rect 950 2174 960 2181
rect 1134 2180 1140 2214
rect 1130 2174 1140 2180
rect 950 2142 1140 2174
rect 950 2108 956 2142
rect 990 2108 1028 2142
rect 1062 2141 1140 2142
rect 1062 2108 1100 2141
rect 950 2107 1100 2108
rect 1134 2107 1140 2141
rect 950 2069 1140 2107
rect 950 2035 956 2069
rect 990 2048 1028 2069
rect 1062 2068 1140 2069
rect 1062 2048 1100 2068
rect 950 1996 960 2035
rect 1134 2034 1140 2068
rect 950 1962 956 1996
rect 1130 1995 1140 2034
rect 950 1923 960 1962
rect 1134 1961 1140 1995
rect 950 1889 956 1923
rect 1130 1922 1140 1961
rect 950 1850 960 1889
rect 1134 1888 1140 1922
rect 950 1816 956 1850
rect 1130 1849 1140 1888
rect 950 1777 960 1816
rect 1134 1815 1140 1849
rect 950 1743 956 1777
rect 1130 1776 1140 1815
rect 950 1704 960 1743
rect 1134 1742 1140 1776
rect 1062 1709 1140 1742
rect 25862 7501 25930 7535
rect 25862 7479 25879 7501
rect 25913 7479 25930 7501
rect 26032 7499 26063 7539
rect 26057 7465 26063 7499
rect 26032 7425 26063 7465
rect 26057 7391 26063 7425
rect 26032 7351 26063 7391
rect 26057 7317 26063 7351
rect 26032 7277 26063 7317
rect 26057 7243 26063 7277
rect 26032 7204 26063 7243
rect 26057 7170 26063 7204
rect 26032 7131 26063 7170
rect 26057 7097 26063 7131
rect 26032 7021 26063 7097
rect 26057 6987 26063 7021
rect 26032 6948 26063 6987
rect 26057 6914 26063 6948
rect 26032 6875 26063 6914
rect 26057 6841 26063 6875
rect 26032 6802 26063 6841
rect 26057 6768 26063 6802
rect 26032 6729 26063 6768
rect 26057 6695 26063 6729
rect 26032 6656 26063 6695
rect 26057 6622 26063 6656
rect 26032 6583 26063 6622
rect 26057 6549 26063 6583
rect 26032 6510 26063 6549
rect 26057 6476 26063 6510
rect 26032 6437 26063 6476
rect 26057 6403 26063 6437
rect 26032 6364 26063 6403
rect 26057 6330 26063 6364
rect 26032 6291 26063 6330
rect 26057 6257 26063 6291
rect 26032 6218 26063 6257
rect 26057 6184 26063 6218
rect 26032 6145 26063 6184
rect 26057 6111 26063 6145
rect 26032 6072 26063 6111
rect 26057 6038 26063 6072
rect 26032 5999 26063 6038
rect 26057 5965 26063 5999
rect 26032 5926 26063 5965
rect 26057 5892 26063 5926
rect 26032 5853 26063 5892
rect 26057 5819 26063 5853
rect 26032 5780 26063 5819
rect 26057 5746 26063 5780
rect 26032 5707 26063 5746
rect 26057 5673 26063 5707
rect 26032 5634 26063 5673
rect 26057 5600 26063 5634
rect 26032 5561 26063 5600
rect 26057 5527 26063 5561
rect 26032 5488 26063 5527
rect 26057 5454 26063 5488
rect 26032 5415 26063 5454
rect 26057 5381 26063 5415
rect 26032 5342 26063 5381
rect 26057 5308 26063 5342
rect 26032 5269 26063 5308
rect 26057 5235 26063 5269
rect 26032 5196 26063 5235
rect 26057 5162 26063 5196
rect 26032 5123 26063 5162
rect 26057 5089 26063 5123
rect 26032 5050 26063 5089
rect 26057 5016 26063 5050
rect 26032 4977 26063 5016
rect 26057 4943 26063 4977
rect 26032 4904 26063 4943
rect 26057 4870 26063 4904
rect 26032 4831 26063 4870
rect 26057 4797 26063 4831
rect 26032 4758 26063 4797
rect 26057 4724 26063 4758
rect 26032 4685 26063 4724
rect 26057 4651 26063 4685
rect 26032 4612 26063 4651
rect 26057 4578 26063 4612
rect 26032 4539 26063 4578
rect 26057 4505 26063 4539
rect 26032 4466 26063 4505
rect 26057 4432 26063 4466
rect 26032 4393 26063 4432
rect 26057 4359 26063 4393
rect 26032 4320 26063 4359
rect 26057 4286 26063 4320
rect 26032 4247 26063 4286
rect 26057 4213 26063 4247
rect 26032 4174 26063 4213
rect 26057 4140 26063 4174
rect 26032 4101 26063 4140
rect 26057 4067 26063 4101
rect 26032 4028 26063 4067
rect 26057 3994 26063 4028
rect 26032 3955 26063 3994
rect 26057 3921 26063 3955
rect 26032 3882 26063 3921
rect 26057 3848 26063 3882
rect 26032 3809 26063 3848
rect 26057 3775 26063 3809
rect 26032 3736 26063 3775
rect 26057 3702 26063 3736
rect 26032 3663 26063 3702
rect 26057 3629 26063 3663
rect 26032 3590 26063 3629
rect 26057 3556 26063 3590
rect 26032 3517 26063 3556
rect 26057 3483 26063 3517
rect 26032 3444 26063 3483
rect 26057 3410 26063 3444
rect 26032 3371 26063 3410
rect 26057 3337 26063 3371
rect 26032 3298 26063 3337
rect 26057 3264 26063 3298
rect 26032 3225 26063 3264
rect 26057 3191 26063 3225
rect 26032 3152 26063 3191
rect 26057 3118 26063 3152
rect 26032 3079 26063 3118
rect 26057 3045 26063 3079
rect 26032 3006 26063 3045
rect 26057 2972 26063 3006
rect 26032 2933 26063 2972
rect 26057 2899 26063 2933
rect 26032 2860 26063 2899
rect 26057 2826 26063 2860
rect 26032 2787 26063 2826
rect 26057 2753 26063 2787
rect 26032 2714 26063 2753
rect 26057 2680 26063 2714
rect 26032 2641 26063 2680
rect 26057 2607 26063 2641
rect 26032 2568 26063 2607
rect 26057 2534 26063 2568
rect 26032 2495 26063 2534
rect 950 1670 956 1704
rect 1062 1703 25862 1709
rect 1062 1699 1100 1703
rect 25110 1699 25149 1703
rect 25183 1699 25222 1703
rect 25256 1699 25295 1703
rect 25329 1699 25368 1703
rect 25402 1699 25441 1703
rect 25475 1699 25514 1703
rect 25548 1699 25587 1703
rect 25621 1699 25660 1703
rect 25694 1699 25733 1703
rect 25767 1699 25806 1703
rect 990 1670 1028 1674
rect 1062 1670 1096 1699
rect 950 1640 1096 1670
rect 950 1631 960 1640
rect 994 1631 1096 1640
rect 25840 1669 25862 1703
rect 25814 1665 25862 1669
rect 25814 1631 25930 1665
rect 950 1597 956 1631
rect 994 1606 1028 1631
rect 990 1597 1028 1606
rect 950 1525 1028 1597
rect 25912 1597 25930 1631
rect 26057 1597 26063 2495
rect 25882 1563 26063 1597
rect 25882 1559 25916 1563
rect 25912 1529 25916 1559
rect 25950 1559 26063 1563
rect 25950 1529 25951 1559
rect 25182 1525 25221 1529
rect 25255 1525 25294 1529
rect 25328 1525 25367 1529
rect 25401 1525 25440 1529
rect 25474 1525 25513 1529
rect 25547 1525 25586 1529
rect 25620 1525 25659 1529
rect 25693 1525 25732 1529
rect 25766 1525 25805 1529
rect 25839 1525 25878 1529
rect 25912 1525 25951 1529
rect 25985 1525 26063 1559
rect 950 1519 26063 1525
rect 26271 7705 26277 7739
rect 26451 7737 26461 7777
rect 26271 7665 26281 7705
rect 26455 7703 26461 7737
rect 26271 7631 26277 7665
rect 26451 7663 26461 7703
rect 26271 7591 26281 7631
rect 26455 7629 26461 7663
rect 26271 7557 26277 7591
rect 26451 7590 26461 7629
rect 26271 7517 26281 7557
rect 26455 7556 26461 7590
rect 26451 7517 26461 7556
rect 26271 7483 26277 7517
rect 26455 7483 26461 7517
rect 26271 7407 26281 7483
rect 26451 7407 26461 7483
rect 26271 7373 26277 7407
rect 26455 7373 26461 7407
rect 26271 7334 26281 7373
rect 26451 7334 26461 7373
rect 26271 7300 26277 7334
rect 26455 7300 26461 7334
rect 26271 7261 26281 7300
rect 26451 7261 26461 7300
rect 26271 7227 26277 7261
rect 26455 7227 26461 7261
rect 26271 7188 26281 7227
rect 26451 7188 26461 7227
rect 26271 7154 26277 7188
rect 26455 7154 26461 7188
rect 26271 7115 26281 7154
rect 26451 7115 26461 7154
rect 26271 7081 26277 7115
rect 26455 7081 26461 7115
rect 26271 7042 26281 7081
rect 26451 7042 26461 7081
rect 564 1437 574 1476
rect 748 1475 754 1509
rect 564 1403 570 1437
rect 744 1436 754 1475
rect 564 1364 574 1403
rect 748 1402 754 1436
rect 564 1330 570 1364
rect 744 1363 754 1402
rect 564 1291 574 1330
rect 748 1329 754 1363
rect 564 1257 570 1291
rect 744 1290 754 1329
rect 564 1218 574 1257
rect 748 1256 754 1290
rect 564 1184 570 1218
rect 744 1217 754 1256
rect 564 1145 574 1184
rect 748 1183 754 1217
rect 564 1111 570 1145
rect 744 1144 754 1183
rect 564 1072 574 1111
rect 748 1110 754 1144
rect 564 1038 570 1072
rect 744 1071 754 1110
rect 564 999 574 1038
rect 748 1037 754 1071
rect 564 965 570 999
rect 744 998 754 1037
rect 564 926 574 965
rect 748 964 754 998
rect 564 892 570 926
rect 744 925 754 964
rect 564 853 574 892
rect 748 891 754 925
rect 564 819 570 853
rect 744 852 754 891
rect 564 780 574 819
rect 748 818 754 852
rect 564 746 570 780
rect 744 779 754 818
rect 564 707 574 746
rect 748 745 754 779
rect 744 730 754 745
rect 26271 730 26277 7042
rect 564 673 570 707
rect 744 706 779 730
rect 813 706 848 730
rect 882 706 917 730
rect 564 634 574 673
rect 676 662 714 696
rect 26315 662 26349 672
rect 676 634 711 662
rect 564 600 570 634
rect 604 600 642 628
rect 564 528 642 600
rect 26455 600 26461 7042
rect 26164 528 26203 560
rect 26237 528 26276 560
rect 26310 528 26349 560
rect 26383 528 26461 600
rect 564 522 26461 528
rect 26674 8099 26680 8133
rect 26858 8099 26864 8133
rect 26674 8054 26684 8099
rect 26854 8054 26864 8099
rect 26674 8020 26680 8054
rect 26858 8020 26864 8054
rect 26674 7975 26684 8020
rect 26854 7975 26864 8020
rect 26674 7941 26680 7975
rect 26858 7941 26864 7975
rect 26674 7896 26684 7941
rect 26854 7896 26864 7941
rect 26674 7862 26680 7896
rect 26858 7862 26864 7896
rect 26674 7786 26684 7862
rect 26854 7786 26864 7862
rect 26674 7752 26680 7786
rect 26858 7752 26864 7786
rect 26674 7713 26684 7752
rect 26854 7713 26864 7752
rect 26674 7679 26680 7713
rect 26858 7679 26864 7713
rect 26674 7640 26684 7679
rect 26854 7640 26864 7679
rect 26674 7606 26680 7640
rect 26858 7606 26864 7640
rect 26674 7567 26684 7606
rect 26854 7567 26864 7606
rect 26674 7533 26680 7567
rect 26858 7533 26864 7567
rect 26674 7494 26684 7533
rect 26854 7494 26864 7533
rect 116 447 122 481
rect 296 480 306 519
rect 116 408 126 447
rect 300 446 306 480
rect 116 374 122 408
rect 296 407 306 446
rect 116 335 126 374
rect 300 373 306 407
rect 296 340 306 373
rect 26674 340 26680 7494
rect 116 301 122 335
rect 296 334 26680 340
rect 116 262 126 301
rect 116 228 122 262
rect 22548 300 22587 334
rect 22621 300 22660 334
rect 22694 300 22733 334
rect 22767 300 22806 334
rect 22840 300 22879 334
rect 22913 300 22952 334
rect 22986 300 23025 334
rect 23059 300 23098 334
rect 23132 300 23171 334
rect 23205 300 23244 334
rect 23278 300 23317 334
rect 23351 300 23390 334
rect 23424 300 23463 334
rect 23497 300 23536 334
rect 23570 300 23609 334
rect 23643 300 23682 334
rect 23716 300 23755 334
rect 23789 300 23828 334
rect 23862 300 23901 334
rect 23935 300 23974 334
rect 24008 300 24047 334
rect 24081 300 24120 334
rect 24154 300 24193 334
rect 24227 300 24266 334
rect 24300 300 24339 334
rect 24373 300 24412 334
rect 24446 300 24485 334
rect 24519 300 24558 334
rect 24592 300 24631 334
rect 24665 300 24704 334
rect 24738 300 24777 334
rect 24811 300 24850 334
rect 24884 300 24923 334
rect 24957 300 24996 334
rect 25030 300 25069 334
rect 25103 300 25142 334
rect 25176 300 25215 334
rect 25249 300 25288 334
rect 25322 300 25361 334
rect 25395 300 25434 334
rect 25468 300 25507 334
rect 25541 300 25580 334
rect 25614 300 25653 334
rect 25687 300 25726 334
rect 25760 300 25799 334
rect 25833 300 25872 334
rect 25906 300 25945 334
rect 25979 300 26018 334
rect 26052 300 26091 334
rect 26125 300 26164 334
rect 26198 300 26237 334
rect 26271 300 26310 334
rect 26344 300 26383 334
rect 26417 300 26456 334
rect 26490 300 26529 334
rect 26563 300 26602 334
rect 26636 300 26680 334
rect 22548 262 26680 300
rect 22548 236 22587 262
rect 22621 236 22660 262
rect 22694 236 22733 262
rect 22767 236 22806 262
rect 22840 236 22879 262
rect 22913 236 22952 262
rect 22986 236 23025 262
rect 23059 236 23098 262
rect 23132 236 23171 262
rect 23205 236 23244 262
rect 23278 236 23317 262
rect 23351 236 23390 262
rect 23424 236 23463 262
rect 23497 236 23536 262
rect 23570 236 23609 262
rect 23643 236 23682 262
rect 23716 236 23755 262
rect 23789 236 23828 262
rect 23862 236 23901 262
rect 23935 236 23974 262
rect 24008 236 24047 262
rect 24081 236 24120 262
rect 24154 236 24193 262
rect 24227 236 24266 262
rect 24300 236 24339 262
rect 24373 236 24412 262
rect 24446 236 24485 262
rect 24519 236 24558 262
rect 24592 236 24631 262
rect 24665 236 24704 262
rect 24738 236 24777 262
rect 24811 236 24850 262
rect 24884 236 24923 262
rect 24957 236 24996 262
rect 25030 236 25069 262
rect 25103 236 25142 262
rect 25176 236 25215 262
rect 25249 236 25288 262
rect 25322 236 25361 262
rect 25395 236 25434 262
rect 25468 236 25507 262
rect 25541 236 25580 262
rect 25614 236 25653 262
rect 25687 236 25726 262
rect 25760 236 25799 262
rect 25833 236 25872 262
rect 25906 236 25945 262
rect 25979 236 26018 262
rect 26052 236 26091 262
rect 26125 236 26164 262
rect 26198 236 26237 262
rect 26271 236 26310 262
rect 26344 236 26383 262
rect 26417 236 26456 262
rect 26490 236 26529 262
rect 26563 236 26602 262
rect 26636 236 26680 262
rect 116 150 126 228
rect 26858 188 26864 7494
rect 126 134 330 140
rect 364 134 399 156
rect 433 134 468 156
rect 502 134 537 156
rect 571 134 606 156
rect 640 134 675 156
rect 709 134 744 156
rect 778 134 813 156
rect 847 134 882 156
rect 916 134 951 156
rect 985 134 1020 156
rect 1054 134 1089 156
rect 1123 134 1158 156
rect 1192 134 1227 156
rect 1261 134 1296 156
rect 1330 134 1365 156
rect 1399 134 1434 156
rect 1468 134 1503 156
rect 1537 134 1572 156
rect 1606 134 1641 156
rect 1675 134 1710 156
rect 1744 134 1779 156
rect 1813 134 1848 156
rect 1882 134 1917 156
rect 1951 134 1986 156
rect 2020 134 2055 156
rect 2089 134 2124 156
rect 2158 134 2193 156
rect 2227 134 2262 156
rect 2296 134 2331 156
rect 2365 134 2400 156
rect 2434 134 2469 156
rect 2503 134 2538 156
rect 2572 134 2607 156
rect 2641 134 2676 156
rect 2710 134 2745 156
rect 2779 134 2814 156
rect 2848 134 2883 156
rect 2917 134 2952 156
rect 126 100 2952 134
rect 26854 150 26864 188
rect 126 66 330 100
rect 364 66 399 100
rect 433 66 468 100
rect 502 66 537 100
rect 571 66 606 100
rect 640 66 675 100
rect 709 66 744 100
rect 778 66 813 100
rect 847 66 882 100
rect 916 66 951 100
rect 985 66 1020 100
rect 1054 66 1089 100
rect 1123 66 1158 100
rect 1192 66 1227 100
rect 1261 66 1296 100
rect 1330 66 1365 100
rect 1399 66 1434 100
rect 1468 66 1503 100
rect 1537 66 1572 100
rect 1606 66 1641 100
rect 1675 66 1710 100
rect 1744 66 1779 100
rect 1813 66 1848 100
rect 1882 66 1917 100
rect 1951 66 1986 100
rect 2020 66 2055 100
rect 2089 66 2124 100
rect 2158 66 2193 100
rect 2227 66 2262 100
rect 2296 66 2331 100
rect 2365 66 2400 100
rect 2434 66 2469 100
rect 2503 66 2538 100
rect 2572 66 2607 100
rect 2641 66 2676 100
rect 2710 66 2745 100
rect 2779 66 2814 100
rect 2848 66 2883 100
rect 2917 66 2952 100
rect 26650 66 26854 100
<< viali >>
rect 194 8470 228 8484
rect 194 8450 228 8470
rect 267 8450 301 8484
rect 340 8450 374 8484
rect 413 8450 447 8484
rect 486 8450 520 8484
rect 559 8450 593 8484
rect 632 8450 666 8484
rect 705 8450 739 8484
rect 778 8450 812 8484
rect 851 8450 885 8484
rect 924 8450 958 8484
rect 997 8450 1031 8484
rect 1070 8450 1104 8484
rect 1143 8450 1177 8484
rect 1216 8450 1250 8484
rect 1289 8450 1323 8484
rect 1362 8450 1396 8484
rect 1435 8450 1469 8484
rect 1508 8450 1542 8484
rect 1581 8450 1615 8484
rect 1654 8450 1688 8484
rect 1727 8450 1761 8484
rect 1800 8450 1834 8484
rect 1873 8450 1907 8484
rect 1946 8450 1980 8484
rect 2019 8450 2053 8484
rect 2092 8450 2126 8484
rect 2165 8450 2199 8484
rect 2238 8450 2272 8484
rect 2311 8450 2345 8484
rect 2384 8450 2418 8484
rect 2457 8450 2491 8484
rect 2530 8450 2564 8484
rect 2603 8450 2637 8484
rect 2676 8450 2710 8484
rect 2749 8450 2783 8484
rect 2822 8450 2856 8484
rect 2895 8450 2929 8484
rect 2968 8450 3002 8484
rect 3041 8450 3075 8484
rect 3114 8450 3148 8484
rect 3187 8450 3221 8484
rect 3260 8450 3294 8484
rect 3333 8450 3367 8484
rect 3406 8450 3440 8484
rect 3479 8450 3513 8484
rect 3552 8450 3586 8484
rect 3625 8450 3659 8484
rect 3698 8450 3732 8484
rect 3771 8450 3805 8484
rect 3844 8450 3878 8484
rect 3917 8450 3951 8484
rect 3990 8450 4024 8484
rect 4063 8450 4097 8484
rect 4136 8450 4170 8484
rect 4209 8450 4243 8484
rect 122 1250 126 8412
rect 126 8340 228 8412
rect 267 8402 301 8412
rect 267 8378 296 8402
rect 296 8378 301 8402
rect 340 8378 374 8412
rect 413 8378 447 8412
rect 486 8378 520 8412
rect 559 8378 593 8412
rect 632 8378 666 8412
rect 705 8378 739 8412
rect 778 8378 812 8412
rect 851 8378 885 8412
rect 924 8378 958 8412
rect 997 8378 1031 8412
rect 1070 8378 1104 8412
rect 1143 8378 1177 8412
rect 1216 8378 1250 8412
rect 1289 8378 1323 8412
rect 1362 8378 1396 8412
rect 1435 8378 1469 8412
rect 1508 8378 1542 8412
rect 1581 8378 1615 8412
rect 1654 8378 1688 8412
rect 1727 8378 1761 8412
rect 1800 8378 1834 8412
rect 1873 8378 1907 8412
rect 1946 8378 1980 8412
rect 2019 8378 2053 8412
rect 2092 8378 2126 8412
rect 2165 8378 2199 8412
rect 2238 8378 2272 8412
rect 2311 8378 2345 8412
rect 2384 8378 2418 8412
rect 2457 8378 2491 8412
rect 2530 8378 2564 8412
rect 2603 8378 2637 8412
rect 2676 8378 2710 8412
rect 2749 8378 2783 8412
rect 2822 8378 2856 8412
rect 2895 8378 2929 8412
rect 2968 8378 3002 8412
rect 3041 8378 3075 8412
rect 3114 8378 3148 8412
rect 3187 8378 3221 8412
rect 3260 8378 3294 8412
rect 3333 8378 3367 8412
rect 3406 8378 3440 8412
rect 3479 8378 3513 8412
rect 3552 8378 3586 8412
rect 3625 8378 3659 8412
rect 3698 8378 3732 8412
rect 3771 8378 3805 8412
rect 3844 8378 3878 8412
rect 3917 8378 3951 8412
rect 3990 8378 4024 8412
rect 4063 8378 4097 8412
rect 4136 8378 4170 8412
rect 4209 8378 4243 8412
rect 4282 8378 26636 8484
rect 26680 8418 26714 8452
rect 26752 8418 26786 8452
rect 26824 8418 26858 8452
rect 4354 8368 26636 8378
rect 26680 8368 26714 8372
rect 126 1322 296 8340
rect 296 1322 300 8340
rect 339 8306 373 8340
rect 412 8306 446 8340
rect 485 8306 519 8340
rect 558 8306 592 8340
rect 631 8306 665 8340
rect 704 8306 738 8340
rect 777 8306 811 8340
rect 850 8306 884 8340
rect 923 8306 957 8340
rect 996 8306 1030 8340
rect 1069 8306 1103 8340
rect 1142 8306 1176 8340
rect 1215 8306 1249 8340
rect 1288 8306 1322 8340
rect 1361 8306 1395 8340
rect 1434 8306 1468 8340
rect 1507 8306 1541 8340
rect 1580 8306 1614 8340
rect 1653 8306 1687 8340
rect 1726 8306 1760 8340
rect 1799 8306 1833 8340
rect 1872 8306 1906 8340
rect 1945 8306 1979 8340
rect 2018 8306 2052 8340
rect 2091 8306 2125 8340
rect 2164 8306 2198 8340
rect 2237 8306 2271 8340
rect 2310 8306 2344 8340
rect 2383 8306 2417 8340
rect 2456 8306 2490 8340
rect 2529 8306 2563 8340
rect 2602 8306 2636 8340
rect 2675 8306 2709 8340
rect 2748 8306 2782 8340
rect 2821 8306 2855 8340
rect 2894 8306 2928 8340
rect 2967 8306 3001 8340
rect 3040 8306 3074 8340
rect 3113 8306 3147 8340
rect 3186 8306 3220 8340
rect 3259 8306 3293 8340
rect 3332 8306 3366 8340
rect 3405 8306 3439 8340
rect 3478 8306 3512 8340
rect 3551 8306 3585 8340
rect 3624 8306 3658 8340
rect 3697 8306 3731 8340
rect 3770 8306 3804 8340
rect 3843 8306 3877 8340
rect 3916 8306 3950 8340
rect 3989 8306 4023 8340
rect 4062 8306 4096 8340
rect 4135 8306 4169 8340
rect 4208 8306 4242 8340
rect 4281 8306 4315 8340
rect 4354 8306 26636 8368
rect 26680 8338 26714 8368
rect 26752 8338 26786 8372
rect 26824 8338 26858 8372
rect 26680 8258 26684 8292
rect 26684 8258 26714 8292
rect 26752 8258 26786 8292
rect 26824 8258 26854 8292
rect 26854 8258 26858 8292
rect 26680 8178 26684 8212
rect 26684 8178 26714 8212
rect 26752 8178 26786 8212
rect 26824 8178 26854 8212
rect 26854 8178 26858 8212
rect 126 1250 228 1322
rect 266 1249 296 1283
rect 296 1249 300 1283
rect 122 1177 126 1211
rect 126 1177 156 1211
rect 194 1177 228 1211
rect 266 1176 296 1210
rect 296 1176 300 1210
rect 122 1104 126 1138
rect 126 1104 156 1138
rect 194 1104 228 1138
rect 266 1103 296 1137
rect 296 1103 300 1137
rect 122 1031 126 1065
rect 126 1031 156 1065
rect 194 1031 228 1065
rect 266 1030 296 1064
rect 296 1030 300 1064
rect 122 958 126 992
rect 126 958 156 992
rect 194 958 228 992
rect 266 957 296 991
rect 296 957 300 991
rect 122 885 126 919
rect 126 885 156 919
rect 194 885 228 919
rect 266 884 296 918
rect 296 884 300 918
rect 122 812 126 846
rect 126 812 156 846
rect 194 812 228 846
rect 266 811 296 845
rect 296 811 300 845
rect 122 739 126 773
rect 126 739 156 773
rect 194 739 228 773
rect 266 738 296 772
rect 296 738 300 772
rect 122 666 126 700
rect 126 666 156 700
rect 194 666 228 700
rect 266 665 296 699
rect 296 665 300 699
rect 122 593 126 627
rect 126 593 156 627
rect 194 593 228 627
rect 266 592 296 626
rect 296 592 300 626
rect 122 520 126 554
rect 126 520 156 554
rect 194 520 228 554
rect 266 519 296 553
rect 296 519 300 553
rect 642 8101 676 8105
rect 715 8101 749 8105
rect 788 8101 822 8105
rect 861 8101 26383 8105
rect 642 8071 676 8101
rect 715 8071 749 8101
rect 788 8071 822 8101
rect 570 7999 574 8033
rect 574 7999 608 8033
rect 608 7999 642 8033
rect 642 7999 676 8033
rect 715 7999 749 8033
rect 788 7999 822 8033
rect 861 7999 26176 8101
rect 26176 8067 26211 8101
rect 26211 8067 26245 8101
rect 26245 8067 26280 8101
rect 26280 8067 26314 8101
rect 26314 8067 26349 8101
rect 26349 8067 26383 8101
rect 26176 8033 26383 8067
rect 26176 7999 26211 8033
rect 26211 7999 26245 8033
rect 26245 7999 26280 8033
rect 26280 7999 26314 8033
rect 26314 7999 26349 8033
rect 26349 7999 26383 8033
rect 26421 7999 26451 8033
rect 26451 7999 26455 8033
rect 570 7964 676 7999
rect 570 7930 574 7964
rect 574 7930 608 7964
rect 608 7930 642 7964
rect 642 7930 676 7964
rect 676 7931 710 7961
rect 710 7931 748 7961
rect 787 7931 821 7961
rect 860 7931 894 7961
rect 933 7931 26108 7999
rect 26108 7965 26311 7999
rect 26108 7931 26143 7965
rect 26143 7931 26177 7965
rect 26177 7931 26212 7965
rect 26212 7931 26246 7965
rect 26246 7931 26281 7965
rect 676 7930 748 7931
rect 570 7896 748 7930
rect 787 7927 821 7931
rect 860 7927 894 7931
rect 933 7927 26281 7931
rect 26281 7927 26311 7965
rect 26349 7925 26383 7959
rect 26421 7925 26451 7959
rect 26451 7925 26455 7959
rect 570 7895 710 7896
rect 570 7861 574 7895
rect 574 7861 608 7895
rect 608 7861 642 7895
rect 642 7861 676 7895
rect 676 7862 710 7895
rect 710 7862 744 7896
rect 744 7862 748 7896
rect 676 7861 748 7862
rect 570 7827 748 7861
rect 570 7826 710 7827
rect 570 7792 574 7826
rect 574 7792 608 7826
rect 608 7792 642 7826
rect 642 7792 676 7826
rect 676 7793 710 7826
rect 710 7793 744 7827
rect 744 7793 748 7827
rect 676 7792 748 7793
rect 570 7758 748 7792
rect 570 7757 710 7758
rect 570 7723 574 7757
rect 574 7723 608 7757
rect 608 7723 642 7757
rect 642 7723 676 7757
rect 676 7724 710 7757
rect 710 7724 744 7758
rect 744 7724 748 7758
rect 676 7723 748 7724
rect 570 7689 748 7723
rect 570 7688 710 7689
rect 570 7654 574 7688
rect 574 7654 608 7688
rect 608 7654 642 7688
rect 642 7654 676 7688
rect 676 7655 710 7688
rect 710 7655 744 7689
rect 744 7655 748 7689
rect 676 7654 748 7655
rect 570 7620 748 7654
rect 570 7619 710 7620
rect 570 7585 574 7619
rect 574 7585 608 7619
rect 608 7585 642 7619
rect 642 7585 676 7619
rect 676 7586 710 7619
rect 710 7586 744 7620
rect 744 7586 748 7620
rect 676 7585 748 7586
rect 570 7551 748 7585
rect 570 7550 710 7551
rect 570 7516 574 7550
rect 574 7516 608 7550
rect 608 7516 642 7550
rect 642 7516 676 7550
rect 676 7517 710 7550
rect 710 7517 744 7551
rect 744 7517 748 7551
rect 676 7516 748 7517
rect 570 7482 748 7516
rect 570 7481 710 7482
rect 570 7447 574 7481
rect 574 7447 608 7481
rect 608 7447 642 7481
rect 642 7447 676 7481
rect 676 7448 710 7481
rect 710 7448 744 7482
rect 744 7448 748 7482
rect 676 7447 748 7448
rect 570 7413 748 7447
rect 570 7412 710 7413
rect 570 7378 574 7412
rect 574 7378 608 7412
rect 608 7378 642 7412
rect 642 7378 676 7412
rect 676 7379 710 7412
rect 710 7379 744 7413
rect 744 7379 748 7413
rect 676 7378 748 7379
rect 570 7344 748 7378
rect 570 7343 710 7344
rect 570 7309 574 7343
rect 574 7309 608 7343
rect 608 7309 642 7343
rect 642 7309 676 7343
rect 676 7310 710 7343
rect 710 7310 744 7344
rect 744 7310 748 7344
rect 676 7309 748 7310
rect 570 7275 748 7309
rect 570 7274 710 7275
rect 570 7240 574 7274
rect 574 7240 608 7274
rect 608 7240 642 7274
rect 642 7240 676 7274
rect 676 7241 710 7274
rect 710 7241 744 7275
rect 744 7241 748 7275
rect 676 7240 748 7241
rect 570 7206 748 7240
rect 570 7205 710 7206
rect 570 7171 574 7205
rect 574 7171 608 7205
rect 608 7171 642 7205
rect 642 7171 676 7205
rect 676 7172 710 7205
rect 710 7172 744 7206
rect 744 7172 748 7206
rect 676 7171 748 7172
rect 570 7137 748 7171
rect 570 7136 710 7137
rect 570 7102 574 7136
rect 574 7102 608 7136
rect 608 7102 642 7136
rect 642 7102 676 7136
rect 676 7103 710 7136
rect 710 7103 744 7137
rect 744 7103 748 7137
rect 676 7102 748 7103
rect 570 7068 748 7102
rect 570 7067 710 7068
rect 570 7033 574 7067
rect 574 7033 608 7067
rect 608 7033 642 7067
rect 642 7033 676 7067
rect 676 7034 710 7067
rect 710 7034 744 7068
rect 744 7034 748 7068
rect 676 7033 748 7034
rect 570 6999 748 7033
rect 570 6998 710 6999
rect 570 6964 574 6998
rect 574 6964 608 6998
rect 608 6964 642 6998
rect 642 6964 676 6998
rect 676 6965 710 6998
rect 710 6965 744 6999
rect 744 6965 748 6999
rect 676 6964 748 6965
rect 570 6930 748 6964
rect 570 6929 710 6930
rect 570 6895 574 6929
rect 574 6895 608 6929
rect 608 6895 642 6929
rect 642 6895 676 6929
rect 676 6896 710 6929
rect 710 6896 744 6930
rect 744 6896 748 6930
rect 676 6895 748 6896
rect 570 6861 748 6895
rect 570 6860 710 6861
rect 570 6826 574 6860
rect 574 6826 608 6860
rect 608 6826 642 6860
rect 642 6826 676 6860
rect 676 6827 710 6860
rect 710 6827 744 6861
rect 744 6827 748 6861
rect 676 6826 748 6827
rect 570 6792 748 6826
rect 570 6791 710 6792
rect 570 6757 574 6791
rect 574 6757 608 6791
rect 608 6757 642 6791
rect 642 6757 676 6791
rect 676 6758 710 6791
rect 710 6758 744 6792
rect 744 6758 748 6792
rect 676 6757 748 6758
rect 570 6723 748 6757
rect 570 6722 710 6723
rect 570 6688 574 6722
rect 574 6688 608 6722
rect 608 6688 642 6722
rect 642 6688 676 6722
rect 676 6689 710 6722
rect 710 6689 744 6723
rect 744 6689 748 6723
rect 676 6688 748 6689
rect 570 6654 748 6688
rect 570 6653 710 6654
rect 570 6619 574 6653
rect 574 6619 608 6653
rect 608 6619 642 6653
rect 642 6619 676 6653
rect 676 6620 710 6653
rect 710 6620 744 6654
rect 744 6620 748 6654
rect 676 6619 748 6620
rect 570 6585 748 6619
rect 570 6584 710 6585
rect 570 6550 574 6584
rect 574 6550 608 6584
rect 608 6550 642 6584
rect 642 6550 676 6584
rect 676 6551 710 6584
rect 710 6551 744 6585
rect 744 6551 748 6585
rect 676 6550 748 6551
rect 570 6516 748 6550
rect 570 6515 710 6516
rect 570 6481 574 6515
rect 574 6481 608 6515
rect 608 6481 642 6515
rect 642 6481 676 6515
rect 676 6482 710 6515
rect 710 6482 744 6516
rect 744 6482 748 6516
rect 676 6481 748 6482
rect 570 6447 748 6481
rect 570 6446 710 6447
rect 570 6412 574 6446
rect 574 6412 608 6446
rect 608 6412 642 6446
rect 642 6412 676 6446
rect 676 6413 710 6446
rect 710 6413 744 6447
rect 744 6413 748 6447
rect 676 6412 748 6413
rect 570 6378 748 6412
rect 570 6377 710 6378
rect 570 6343 574 6377
rect 574 6343 608 6377
rect 608 6343 642 6377
rect 642 6343 676 6377
rect 676 6344 710 6377
rect 710 6344 744 6378
rect 744 6344 748 6378
rect 676 6343 748 6344
rect 570 6309 748 6343
rect 570 6308 710 6309
rect 570 6274 574 6308
rect 574 6274 608 6308
rect 608 6274 642 6308
rect 642 6274 676 6308
rect 676 6275 710 6308
rect 710 6275 744 6309
rect 744 6275 748 6309
rect 676 6274 748 6275
rect 570 6240 748 6274
rect 570 6239 710 6240
rect 570 6205 574 6239
rect 574 6205 608 6239
rect 608 6205 642 6239
rect 642 6205 676 6239
rect 676 6206 710 6239
rect 710 6206 744 6240
rect 744 6206 748 6240
rect 676 6205 748 6206
rect 570 6171 748 6205
rect 570 6170 710 6171
rect 570 6136 574 6170
rect 574 6136 608 6170
rect 608 6136 642 6170
rect 642 6136 676 6170
rect 676 6137 710 6170
rect 710 6137 744 6171
rect 744 6137 748 6171
rect 676 6136 748 6137
rect 570 6102 748 6136
rect 570 6101 710 6102
rect 570 6067 574 6101
rect 574 6067 608 6101
rect 608 6067 642 6101
rect 642 6067 676 6101
rect 676 6068 710 6101
rect 710 6068 744 6102
rect 744 6068 748 6102
rect 676 6067 748 6068
rect 570 6033 748 6067
rect 570 6032 710 6033
rect 570 5998 574 6032
rect 574 5998 608 6032
rect 608 5998 642 6032
rect 642 5998 676 6032
rect 676 5999 710 6032
rect 710 5999 744 6033
rect 744 5999 748 6033
rect 676 5998 748 5999
rect 570 5964 748 5998
rect 570 5963 710 5964
rect 570 5929 574 5963
rect 574 5929 608 5963
rect 608 5929 642 5963
rect 642 5929 676 5963
rect 676 5930 710 5963
rect 710 5930 744 5964
rect 744 5930 748 5964
rect 676 5929 748 5930
rect 570 5895 748 5929
rect 570 5894 710 5895
rect 570 5860 574 5894
rect 574 5860 608 5894
rect 608 5860 642 5894
rect 642 5860 676 5894
rect 676 5861 710 5894
rect 710 5861 744 5895
rect 744 5861 748 5895
rect 676 5860 748 5861
rect 570 5826 748 5860
rect 570 5825 710 5826
rect 570 5791 574 5825
rect 574 5791 608 5825
rect 608 5791 642 5825
rect 642 5791 676 5825
rect 676 5792 710 5825
rect 710 5792 744 5826
rect 744 5792 748 5826
rect 676 5791 748 5792
rect 570 5757 748 5791
rect 570 5756 710 5757
rect 570 5722 574 5756
rect 574 5722 608 5756
rect 608 5722 642 5756
rect 642 5722 676 5756
rect 676 5723 710 5756
rect 710 5723 744 5757
rect 744 5723 748 5757
rect 676 5722 748 5723
rect 570 5688 748 5722
rect 570 5687 710 5688
rect 570 5653 574 5687
rect 574 5653 608 5687
rect 608 5653 642 5687
rect 642 5653 676 5687
rect 676 5654 710 5687
rect 710 5654 744 5688
rect 744 5654 748 5688
rect 676 5653 748 5654
rect 570 5619 748 5653
rect 570 5618 710 5619
rect 570 5584 574 5618
rect 574 5584 608 5618
rect 608 5584 642 5618
rect 642 5584 676 5618
rect 676 5585 710 5618
rect 710 5585 744 5619
rect 744 5585 748 5619
rect 676 5584 748 5585
rect 570 5550 748 5584
rect 570 5549 710 5550
rect 570 5515 574 5549
rect 574 5515 608 5549
rect 608 5515 642 5549
rect 642 5515 676 5549
rect 676 5516 710 5549
rect 710 5516 744 5550
rect 744 5516 748 5550
rect 676 5515 748 5516
rect 570 5481 748 5515
rect 570 5480 710 5481
rect 570 5446 574 5480
rect 574 5446 608 5480
rect 608 5446 642 5480
rect 642 5446 676 5480
rect 676 5447 710 5480
rect 710 5447 744 5481
rect 744 5447 748 5481
rect 676 5446 748 5447
rect 570 5412 748 5446
rect 570 5411 710 5412
rect 570 5377 574 5411
rect 574 5377 608 5411
rect 608 5377 642 5411
rect 642 5377 676 5411
rect 676 5378 710 5411
rect 710 5378 744 5412
rect 744 5378 748 5412
rect 676 5377 748 5378
rect 570 5343 748 5377
rect 570 5342 710 5343
rect 570 5308 574 5342
rect 574 5308 608 5342
rect 608 5308 642 5342
rect 642 5308 676 5342
rect 676 5309 710 5342
rect 710 5309 744 5343
rect 744 5309 748 5343
rect 676 5308 748 5309
rect 570 5274 748 5308
rect 570 5273 710 5274
rect 570 4695 574 5273
rect 574 5205 676 5273
rect 676 5240 710 5273
rect 710 5240 744 5274
rect 744 5240 748 5274
rect 676 5205 748 5240
rect 574 4695 744 5205
rect 744 4695 748 5205
rect 570 4687 748 4695
rect 26277 7853 26281 7887
rect 26281 7853 26311 7887
rect 26349 7851 26383 7885
rect 26421 7851 26451 7885
rect 26451 7851 26455 7885
rect 26277 7779 26281 7813
rect 26281 7779 26311 7813
rect 26349 7777 26383 7811
rect 26421 7777 26451 7811
rect 26451 7777 26455 7811
rect 570 4627 676 4687
rect 714 4627 748 4648
rect 570 4615 574 4627
rect 574 4615 608 4627
rect 608 4615 642 4627
rect 642 4615 676 4627
rect 714 4614 744 4627
rect 744 4614 748 4627
rect 570 4558 604 4576
rect 642 4558 676 4576
rect 714 4558 748 4575
rect 570 4542 574 4558
rect 574 4542 604 4558
rect 642 4542 676 4558
rect 714 4541 744 4558
rect 744 4541 748 4558
rect 570 4489 604 4503
rect 642 4489 676 4503
rect 714 4489 748 4502
rect 570 4469 574 4489
rect 574 4469 604 4489
rect 642 4469 676 4489
rect 714 4468 744 4489
rect 744 4468 748 4489
rect 570 4420 604 4430
rect 642 4420 676 4430
rect 714 4420 748 4429
rect 570 4396 574 4420
rect 574 4396 604 4420
rect 642 4396 676 4420
rect 714 4395 744 4420
rect 744 4395 748 4420
rect 570 4351 604 4357
rect 642 4351 676 4357
rect 714 4351 748 4356
rect 570 4323 574 4351
rect 574 4323 604 4351
rect 642 4323 676 4351
rect 714 4322 744 4351
rect 744 4322 748 4351
rect 570 4282 604 4284
rect 642 4282 676 4284
rect 714 4282 748 4283
rect 570 4250 574 4282
rect 574 4250 604 4282
rect 642 4250 676 4282
rect 714 4249 744 4282
rect 744 4249 748 4282
rect 570 4179 574 4211
rect 574 4179 604 4211
rect 642 4179 676 4211
rect 714 4179 744 4210
rect 744 4179 748 4210
rect 570 4177 604 4179
rect 642 4177 676 4179
rect 714 4176 748 4179
rect 570 4110 574 4138
rect 574 4110 604 4138
rect 642 4110 676 4138
rect 714 4110 744 4137
rect 744 4110 748 4137
rect 570 4104 604 4110
rect 642 4104 676 4110
rect 714 4103 748 4110
rect 570 4041 574 4065
rect 574 4041 604 4065
rect 642 4041 676 4065
rect 714 4041 744 4064
rect 744 4041 748 4064
rect 570 4031 604 4041
rect 642 4031 676 4041
rect 714 4030 748 4041
rect 570 3972 574 3992
rect 574 3972 604 3992
rect 642 3972 676 3992
rect 714 3972 744 3991
rect 744 3972 748 3991
rect 570 3958 604 3972
rect 642 3958 676 3972
rect 714 3957 748 3972
rect 570 3903 574 3919
rect 574 3903 604 3919
rect 642 3903 676 3919
rect 714 3903 744 3918
rect 744 3903 748 3918
rect 570 3885 604 3903
rect 642 3885 676 3903
rect 714 3884 748 3903
rect 570 3834 574 3846
rect 574 3834 604 3846
rect 642 3834 676 3846
rect 714 3834 744 3845
rect 744 3834 748 3845
rect 570 3812 604 3834
rect 642 3812 676 3834
rect 714 3811 748 3834
rect 570 3765 574 3773
rect 574 3765 604 3773
rect 642 3765 676 3773
rect 714 3765 744 3772
rect 744 3765 748 3772
rect 570 3739 604 3765
rect 642 3739 676 3765
rect 714 3738 748 3765
rect 570 3696 574 3700
rect 574 3696 604 3700
rect 642 3696 676 3700
rect 714 3696 744 3699
rect 744 3696 748 3699
rect 570 3666 604 3696
rect 642 3666 676 3696
rect 714 3665 748 3696
rect 570 3593 604 3627
rect 642 3593 676 3627
rect 714 3592 748 3626
rect 570 3523 604 3554
rect 642 3523 676 3554
rect 714 3523 748 3553
rect 570 3520 574 3523
rect 574 3520 604 3523
rect 642 3520 676 3523
rect 714 3519 744 3523
rect 744 3519 748 3523
rect 570 3454 604 3481
rect 642 3454 676 3481
rect 714 3454 748 3480
rect 570 3447 574 3454
rect 574 3447 604 3454
rect 642 3447 676 3454
rect 714 3446 744 3454
rect 744 3446 748 3454
rect 570 3385 604 3408
rect 642 3385 676 3408
rect 714 3385 748 3407
rect 570 3374 574 3385
rect 574 3374 604 3385
rect 642 3374 676 3385
rect 714 3373 744 3385
rect 744 3373 748 3385
rect 570 3316 604 3335
rect 642 3316 676 3335
rect 714 3316 748 3334
rect 570 3301 574 3316
rect 574 3301 604 3316
rect 642 3301 676 3316
rect 714 3300 744 3316
rect 744 3300 748 3316
rect 570 3247 604 3262
rect 642 3247 676 3262
rect 714 3247 748 3261
rect 570 3228 574 3247
rect 574 3228 604 3247
rect 642 3228 676 3247
rect 714 3227 744 3247
rect 744 3227 748 3247
rect 570 3178 604 3189
rect 642 3178 676 3189
rect 714 3178 748 3188
rect 570 3155 574 3178
rect 574 3155 604 3178
rect 642 3155 676 3178
rect 714 3154 744 3178
rect 744 3154 748 3178
rect 570 3082 574 3116
rect 574 3082 604 3116
rect 642 3082 676 3116
rect 714 3081 744 3115
rect 744 3081 748 3115
rect 570 3009 574 3043
rect 574 3009 604 3043
rect 642 3009 676 3043
rect 714 3008 744 3042
rect 744 3008 748 3042
rect 570 2936 574 2970
rect 574 2936 604 2970
rect 642 2936 676 2970
rect 714 2935 744 2969
rect 744 2935 748 2969
rect 570 2863 574 2897
rect 574 2863 604 2897
rect 642 2863 676 2897
rect 714 2862 744 2896
rect 744 2862 748 2896
rect 570 2790 574 2824
rect 574 2790 604 2824
rect 642 2790 676 2824
rect 714 2789 744 2823
rect 744 2789 748 2823
rect 570 2717 574 2751
rect 574 2717 604 2751
rect 642 2717 676 2751
rect 714 2716 744 2750
rect 744 2716 748 2750
rect 570 2644 574 2678
rect 574 2644 604 2678
rect 642 2644 676 2678
rect 714 2643 744 2677
rect 744 2643 748 2677
rect 570 2571 574 2605
rect 574 2571 604 2605
rect 642 2571 676 2605
rect 714 2570 744 2604
rect 744 2570 748 2604
rect 570 2498 574 2532
rect 574 2498 604 2532
rect 642 2498 676 2532
rect 714 2497 744 2531
rect 744 2497 748 2531
rect 570 2425 574 2459
rect 574 2425 604 2459
rect 642 2425 676 2459
rect 714 2424 744 2458
rect 744 2424 748 2458
rect 570 2352 574 2386
rect 574 2352 604 2386
rect 642 2352 676 2386
rect 714 2351 744 2385
rect 744 2351 748 2385
rect 570 2279 574 2313
rect 574 2279 604 2313
rect 642 2279 676 2313
rect 714 2278 744 2312
rect 744 2278 748 2312
rect 570 2206 574 2240
rect 574 2206 604 2240
rect 642 2206 676 2240
rect 714 2205 744 2239
rect 744 2205 748 2239
rect 570 2133 574 2167
rect 574 2133 604 2167
rect 642 2133 676 2167
rect 714 2132 744 2166
rect 744 2132 748 2166
rect 570 2060 574 2094
rect 574 2060 604 2094
rect 642 2060 676 2094
rect 714 2059 744 2093
rect 744 2059 748 2093
rect 570 1987 574 2021
rect 574 1987 604 2021
rect 642 1987 676 2021
rect 714 1986 744 2020
rect 744 1986 748 2020
rect 570 1914 574 1948
rect 574 1914 604 1948
rect 642 1914 676 1948
rect 714 1913 744 1947
rect 744 1913 748 1947
rect 570 1841 574 1875
rect 574 1841 604 1875
rect 642 1841 676 1875
rect 714 1840 744 1874
rect 744 1840 748 1874
rect 570 1768 574 1802
rect 574 1768 604 1802
rect 642 1768 676 1802
rect 714 1767 744 1801
rect 744 1767 748 1801
rect 570 1695 574 1729
rect 574 1695 604 1729
rect 642 1695 676 1729
rect 714 1694 744 1728
rect 744 1694 748 1728
rect 570 1622 574 1656
rect 574 1622 604 1656
rect 642 1622 676 1656
rect 714 1621 744 1655
rect 744 1621 748 1655
rect 570 1549 574 1583
rect 574 1549 604 1583
rect 642 1549 676 1583
rect 714 1548 744 1582
rect 744 1548 748 1582
rect 570 1476 574 1510
rect 574 1476 604 1510
rect 642 1476 676 1510
rect 1028 7716 1062 7719
rect 1101 7716 1135 7719
rect 1174 7716 1208 7719
rect 1247 7716 1281 7719
rect 1320 7716 1354 7719
rect 1393 7716 1427 7719
rect 1466 7716 1500 7719
rect 1539 7716 1573 7719
rect 1612 7716 1646 7719
rect 1685 7716 1719 7719
rect 1758 7716 1792 7719
rect 1831 7716 25985 7719
rect 1028 7685 1042 7716
rect 1042 7685 1062 7716
rect 1101 7685 1110 7716
rect 1110 7685 1135 7716
rect 1174 7685 1208 7716
rect 1247 7685 1281 7716
rect 1320 7685 1354 7716
rect 1393 7685 1427 7716
rect 1466 7685 1500 7716
rect 1539 7685 1573 7716
rect 1612 7685 1646 7716
rect 1685 7685 1719 7716
rect 1758 7685 1792 7716
rect 956 4517 960 7647
rect 960 7575 1062 7647
rect 1101 7614 1110 7647
rect 1110 7614 1135 7647
rect 1174 7614 1208 7647
rect 1101 7613 1135 7614
rect 1174 7613 1178 7614
rect 1178 7613 1208 7614
rect 1247 7613 1281 7647
rect 1320 7613 1354 7647
rect 1393 7613 1427 7647
rect 1466 7613 1500 7647
rect 1539 7613 1573 7647
rect 1612 7613 1646 7647
rect 1685 7613 1719 7647
rect 1758 7613 1792 7647
rect 1831 7614 25964 7716
rect 25964 7614 25985 7716
rect 26023 7615 26057 7647
rect 1831 7613 25896 7614
rect 25896 7613 25985 7614
rect 26023 7613 26032 7615
rect 26032 7613 26057 7615
rect 960 4589 1130 7575
rect 1130 4589 1134 7575
rect 1173 7546 1178 7575
rect 1178 7546 1207 7575
rect 1246 7546 1280 7575
rect 1319 7546 1353 7575
rect 1392 7546 1426 7575
rect 1465 7546 1499 7575
rect 1538 7546 1572 7575
rect 1611 7546 1645 7575
rect 1684 7546 1718 7575
rect 1757 7546 1791 7575
rect 1830 7546 1864 7575
rect 1903 7546 25896 7613
rect 25896 7546 25913 7613
rect 25951 7547 25985 7573
rect 26023 7547 26057 7573
rect 1173 7541 1207 7546
rect 1246 7541 1280 7546
rect 1319 7541 1353 7546
rect 1392 7541 1426 7546
rect 1465 7541 1499 7546
rect 1538 7541 1572 7546
rect 1611 7541 1645 7546
rect 1684 7541 1718 7546
rect 1757 7541 1791 7546
rect 1830 7541 1864 7546
rect 1903 7541 25913 7546
rect 25951 7539 25985 7547
rect 26023 7539 26032 7547
rect 26032 7539 26057 7547
rect 960 4517 1062 4589
rect 1100 4516 1130 4550
rect 1130 4516 1134 4550
rect 956 4444 960 4478
rect 960 4444 990 4478
rect 1028 4444 1062 4478
rect 1100 4443 1130 4477
rect 1130 4443 1134 4477
rect 956 4371 960 4405
rect 960 4371 990 4405
rect 1028 4371 1062 4405
rect 1100 4370 1130 4404
rect 1130 4370 1134 4404
rect 956 4298 960 4332
rect 960 4298 990 4332
rect 1028 4298 1062 4332
rect 1100 4297 1130 4331
rect 1130 4297 1134 4331
rect 956 4225 960 4259
rect 960 4225 990 4259
rect 1028 4225 1062 4259
rect 1100 4224 1130 4258
rect 1130 4224 1134 4258
rect 956 4152 960 4186
rect 960 4152 990 4186
rect 1028 4152 1062 4186
rect 1100 4151 1130 4185
rect 1130 4151 1134 4185
rect 956 4079 960 4113
rect 960 4079 990 4113
rect 1028 4079 1062 4113
rect 1100 4078 1130 4112
rect 1130 4078 1134 4112
rect 956 4006 960 4040
rect 960 4006 990 4040
rect 1028 4006 1062 4040
rect 1100 4005 1130 4039
rect 1130 4005 1134 4039
rect 956 3933 960 3967
rect 960 3933 990 3967
rect 1028 3933 1062 3967
rect 1100 3932 1130 3966
rect 1130 3932 1134 3966
rect 956 3860 960 3894
rect 960 3860 990 3894
rect 1028 3860 1062 3894
rect 1100 3859 1130 3893
rect 1130 3859 1134 3893
rect 956 3787 960 3821
rect 960 3787 990 3821
rect 1028 3787 1062 3821
rect 1100 3786 1130 3820
rect 1130 3786 1134 3820
rect 956 3714 960 3748
rect 960 3714 990 3748
rect 1028 3714 1062 3748
rect 1100 3713 1130 3747
rect 1130 3713 1134 3747
rect 956 3641 960 3675
rect 960 3641 990 3675
rect 1028 3641 1062 3675
rect 1100 3640 1130 3674
rect 1130 3640 1134 3674
rect 956 3568 960 3602
rect 960 3568 990 3602
rect 1028 3568 1062 3602
rect 1100 3567 1130 3601
rect 1130 3567 1134 3601
rect 956 3495 960 3529
rect 960 3495 990 3529
rect 1028 3495 1062 3529
rect 1100 3494 1130 3528
rect 1130 3494 1134 3528
rect 956 3422 960 3456
rect 960 3422 990 3456
rect 1028 3422 1062 3456
rect 1100 3421 1130 3455
rect 1130 3421 1134 3455
rect 956 3349 960 3383
rect 960 3349 990 3383
rect 1028 3349 1062 3383
rect 1100 3348 1130 3382
rect 1130 3348 1134 3382
rect 956 3276 960 3310
rect 960 3276 990 3310
rect 1028 3276 1062 3310
rect 1100 3275 1130 3309
rect 1130 3275 1134 3309
rect 956 3203 960 3237
rect 960 3203 990 3237
rect 1028 3203 1062 3237
rect 1100 3202 1130 3236
rect 1130 3202 1134 3236
rect 956 3130 960 3164
rect 960 3130 990 3164
rect 1028 3130 1062 3164
rect 1100 3129 1130 3163
rect 1130 3129 1134 3163
rect 956 3057 960 3091
rect 960 3057 990 3091
rect 1028 3057 1062 3091
rect 1100 3056 1130 3090
rect 1130 3056 1134 3090
rect 956 2984 960 3018
rect 960 2984 990 3018
rect 1028 2984 1062 3018
rect 1100 2983 1130 3017
rect 1130 2983 1134 3017
rect 956 2911 960 2945
rect 960 2911 990 2945
rect 1028 2911 1062 2945
rect 1100 2910 1130 2944
rect 1130 2910 1134 2944
rect 956 2838 960 2872
rect 960 2838 990 2872
rect 1028 2838 1062 2872
rect 1100 2837 1130 2871
rect 1130 2837 1134 2871
rect 956 2765 960 2799
rect 960 2765 990 2799
rect 1028 2765 1062 2799
rect 1100 2764 1130 2798
rect 1130 2764 1134 2798
rect 956 2692 960 2726
rect 960 2692 990 2726
rect 1028 2692 1062 2726
rect 1100 2691 1130 2725
rect 1130 2691 1134 2725
rect 956 2619 960 2653
rect 960 2619 990 2653
rect 1028 2619 1062 2653
rect 1100 2618 1130 2652
rect 1130 2618 1134 2652
rect 956 2546 960 2580
rect 960 2546 990 2580
rect 1028 2546 1062 2580
rect 1100 2545 1130 2579
rect 1130 2545 1134 2579
rect 956 2473 960 2507
rect 960 2473 990 2507
rect 1028 2473 1062 2507
rect 1100 2472 1130 2506
rect 1130 2472 1134 2506
rect 956 2400 960 2434
rect 960 2400 990 2434
rect 1028 2400 1062 2434
rect 1100 2399 1130 2433
rect 1130 2399 1134 2433
rect 956 2327 960 2361
rect 960 2327 990 2361
rect 1028 2327 1062 2361
rect 1100 2326 1130 2360
rect 1130 2326 1134 2360
rect 956 2254 960 2288
rect 960 2254 990 2288
rect 1028 2254 1062 2288
rect 1100 2253 1130 2287
rect 1130 2253 1134 2287
rect 956 2181 960 2215
rect 960 2181 990 2215
rect 1028 2181 1062 2215
rect 1100 2180 1130 2214
rect 1130 2180 1134 2214
rect 956 2108 990 2142
rect 1028 2108 1062 2142
rect 1100 2107 1134 2141
rect 956 2048 990 2069
rect 1028 2048 1062 2069
rect 1100 2048 1134 2068
rect 956 2035 960 2048
rect 960 2035 990 2048
rect 1028 2035 1062 2048
rect 1100 2034 1130 2048
rect 1130 2034 1134 2048
rect 956 1962 960 1996
rect 960 1962 990 1996
rect 1028 1962 1062 1996
rect 1100 1961 1130 1995
rect 1130 1961 1134 1995
rect 956 1889 960 1923
rect 960 1889 990 1923
rect 1028 1889 1062 1923
rect 1100 1888 1130 1922
rect 1130 1888 1134 1922
rect 956 1816 960 1850
rect 960 1816 990 1850
rect 1028 1816 1062 1850
rect 1100 1815 1130 1849
rect 1130 1815 1134 1849
rect 956 1743 960 1777
rect 960 1743 990 1777
rect 1028 1743 1062 1777
rect 1100 1742 1130 1776
rect 1130 1742 1134 1776
rect 25879 7479 25913 7501
rect 25879 7467 25913 7479
rect 25951 7465 25985 7499
rect 26023 7465 26032 7499
rect 26032 7465 26057 7499
rect 25879 7393 25913 7427
rect 25951 7391 25985 7425
rect 26023 7391 26032 7425
rect 26032 7391 26057 7425
rect 25879 7319 25913 7353
rect 25951 7317 25985 7351
rect 26023 7317 26032 7351
rect 26032 7317 26057 7351
rect 25879 7245 25913 7279
rect 25951 7243 25985 7277
rect 26023 7243 26032 7277
rect 26032 7243 26057 7277
rect 25879 7171 25913 7205
rect 25951 7170 25985 7204
rect 26023 7170 26032 7204
rect 26032 7170 26057 7204
rect 25879 7097 25913 7131
rect 25951 7097 25985 7131
rect 26023 7097 26032 7131
rect 26032 7097 26057 7131
rect 25879 6987 25913 7021
rect 25951 6987 25985 7021
rect 26023 6987 26032 7021
rect 26032 6987 26057 7021
rect 25879 6914 25913 6948
rect 25951 6914 25985 6948
rect 26023 6914 26032 6948
rect 26032 6914 26057 6948
rect 25879 6841 25913 6875
rect 25951 6841 25985 6875
rect 26023 6841 26032 6875
rect 26032 6841 26057 6875
rect 25879 6768 25913 6802
rect 25951 6768 25985 6802
rect 26023 6768 26032 6802
rect 26032 6768 26057 6802
rect 25879 6695 25913 6729
rect 25951 6695 25985 6729
rect 26023 6695 26032 6729
rect 26032 6695 26057 6729
rect 25879 6622 25913 6656
rect 25951 6622 25985 6656
rect 26023 6622 26032 6656
rect 26032 6622 26057 6656
rect 25879 6549 25913 6583
rect 25951 6549 25985 6583
rect 26023 6549 26032 6583
rect 26032 6549 26057 6583
rect 25879 6476 25913 6510
rect 25951 6476 25985 6510
rect 26023 6476 26032 6510
rect 26032 6476 26057 6510
rect 25879 6403 25913 6437
rect 25951 6403 25985 6437
rect 26023 6403 26032 6437
rect 26032 6403 26057 6437
rect 25879 6330 25913 6364
rect 25951 6330 25985 6364
rect 26023 6330 26032 6364
rect 26032 6330 26057 6364
rect 25879 6257 25913 6291
rect 25951 6257 25985 6291
rect 26023 6257 26032 6291
rect 26032 6257 26057 6291
rect 25879 6184 25913 6218
rect 25951 6184 25985 6218
rect 26023 6184 26032 6218
rect 26032 6184 26057 6218
rect 25879 6111 25913 6145
rect 25951 6111 25985 6145
rect 26023 6111 26032 6145
rect 26032 6111 26057 6145
rect 25879 6038 25913 6072
rect 25951 6038 25985 6072
rect 26023 6038 26032 6072
rect 26032 6038 26057 6072
rect 25879 5965 25913 5999
rect 25951 5965 25985 5999
rect 26023 5965 26032 5999
rect 26032 5965 26057 5999
rect 25879 5892 25913 5926
rect 25951 5892 25985 5926
rect 26023 5892 26032 5926
rect 26032 5892 26057 5926
rect 25879 5819 25913 5853
rect 25951 5819 25985 5853
rect 26023 5819 26032 5853
rect 26032 5819 26057 5853
rect 25879 5746 25913 5780
rect 25951 5746 25985 5780
rect 26023 5746 26032 5780
rect 26032 5746 26057 5780
rect 25879 5673 25913 5707
rect 25951 5673 25985 5707
rect 26023 5673 26032 5707
rect 26032 5673 26057 5707
rect 25879 5600 25913 5634
rect 25951 5600 25985 5634
rect 26023 5600 26032 5634
rect 26032 5600 26057 5634
rect 25879 5527 25913 5561
rect 25951 5527 25985 5561
rect 26023 5527 26032 5561
rect 26032 5527 26057 5561
rect 25879 5454 25913 5488
rect 25951 5454 25985 5488
rect 26023 5454 26032 5488
rect 26032 5454 26057 5488
rect 25879 5381 25913 5415
rect 25951 5381 25985 5415
rect 26023 5381 26032 5415
rect 26032 5381 26057 5415
rect 25879 5308 25913 5342
rect 25951 5308 25985 5342
rect 26023 5308 26032 5342
rect 26032 5308 26057 5342
rect 25879 5235 25913 5269
rect 25951 5235 25985 5269
rect 26023 5235 26032 5269
rect 26032 5235 26057 5269
rect 25879 5162 25913 5196
rect 25951 5162 25985 5196
rect 26023 5162 26032 5196
rect 26032 5162 26057 5196
rect 25879 5089 25913 5123
rect 25951 5089 25985 5123
rect 26023 5089 26032 5123
rect 26032 5089 26057 5123
rect 25879 5016 25913 5050
rect 25951 5016 25985 5050
rect 26023 5016 26032 5050
rect 26032 5016 26057 5050
rect 25879 4943 25913 4977
rect 25951 4943 25985 4977
rect 26023 4943 26032 4977
rect 26032 4943 26057 4977
rect 25879 4870 25913 4904
rect 25951 4870 25985 4904
rect 26023 4870 26032 4904
rect 26032 4870 26057 4904
rect 25879 4797 25913 4831
rect 25951 4797 25985 4831
rect 26023 4797 26032 4831
rect 26032 4797 26057 4831
rect 25879 4724 25913 4758
rect 25951 4724 25985 4758
rect 26023 4724 26032 4758
rect 26032 4724 26057 4758
rect 25879 4651 25913 4685
rect 25951 4651 25985 4685
rect 26023 4651 26032 4685
rect 26032 4651 26057 4685
rect 25879 4578 25913 4612
rect 25951 4578 25985 4612
rect 26023 4578 26032 4612
rect 26032 4578 26057 4612
rect 25879 4505 25913 4539
rect 25951 4505 25985 4539
rect 26023 4505 26032 4539
rect 26032 4505 26057 4539
rect 25879 4432 25913 4466
rect 25951 4432 25985 4466
rect 26023 4432 26032 4466
rect 26032 4432 26057 4466
rect 25879 4359 25913 4393
rect 25951 4359 25985 4393
rect 26023 4359 26032 4393
rect 26032 4359 26057 4393
rect 25879 4286 25913 4320
rect 25951 4286 25985 4320
rect 26023 4286 26032 4320
rect 26032 4286 26057 4320
rect 25879 4213 25913 4247
rect 25951 4213 25985 4247
rect 26023 4213 26032 4247
rect 26032 4213 26057 4247
rect 25879 4140 25913 4174
rect 25951 4140 25985 4174
rect 26023 4140 26032 4174
rect 26032 4140 26057 4174
rect 25879 4067 25913 4101
rect 25951 4067 25985 4101
rect 26023 4067 26032 4101
rect 26032 4067 26057 4101
rect 25879 3994 25913 4028
rect 25951 3994 25985 4028
rect 26023 3994 26032 4028
rect 26032 3994 26057 4028
rect 25879 3921 25913 3955
rect 25951 3921 25985 3955
rect 26023 3921 26032 3955
rect 26032 3921 26057 3955
rect 25879 3848 25913 3882
rect 25951 3848 25985 3882
rect 26023 3848 26032 3882
rect 26032 3848 26057 3882
rect 25879 3775 25913 3809
rect 25951 3775 25985 3809
rect 26023 3775 26032 3809
rect 26032 3775 26057 3809
rect 25879 3702 25913 3736
rect 25951 3702 25985 3736
rect 26023 3702 26032 3736
rect 26032 3702 26057 3736
rect 25879 3629 25913 3663
rect 25951 3629 25985 3663
rect 26023 3629 26032 3663
rect 26032 3629 26057 3663
rect 25879 3556 25913 3590
rect 25951 3556 25985 3590
rect 26023 3556 26032 3590
rect 26032 3556 26057 3590
rect 25879 3483 25913 3517
rect 25951 3483 25985 3517
rect 26023 3483 26032 3517
rect 26032 3483 26057 3517
rect 25879 3410 25913 3444
rect 25951 3410 25985 3444
rect 26023 3410 26032 3444
rect 26032 3410 26057 3444
rect 25879 3337 25913 3371
rect 25951 3337 25985 3371
rect 26023 3337 26032 3371
rect 26032 3337 26057 3371
rect 25879 3264 25913 3298
rect 25951 3264 25985 3298
rect 26023 3264 26032 3298
rect 26032 3264 26057 3298
rect 25879 3191 25913 3225
rect 25951 3191 25985 3225
rect 26023 3191 26032 3225
rect 26032 3191 26057 3225
rect 25879 3118 25913 3152
rect 25951 3118 25985 3152
rect 26023 3118 26032 3152
rect 26032 3118 26057 3152
rect 25879 3045 25913 3079
rect 25951 3045 25985 3079
rect 26023 3045 26032 3079
rect 26032 3045 26057 3079
rect 25879 2972 25913 3006
rect 25951 2972 25985 3006
rect 26023 2972 26032 3006
rect 26032 2972 26057 3006
rect 25879 2899 25913 2933
rect 25951 2899 25985 2933
rect 26023 2899 26032 2933
rect 26032 2899 26057 2933
rect 25879 2826 25913 2860
rect 25951 2826 25985 2860
rect 26023 2826 26032 2860
rect 26032 2826 26057 2860
rect 25879 2753 25913 2787
rect 25951 2753 25985 2787
rect 26023 2753 26032 2787
rect 26032 2753 26057 2787
rect 25879 2680 25913 2714
rect 25951 2680 25985 2714
rect 26023 2680 26032 2714
rect 26032 2680 26057 2714
rect 25879 2607 25913 2641
rect 25951 2607 25985 2641
rect 26023 2607 26032 2641
rect 26032 2607 26057 2641
rect 25879 2534 25913 2568
rect 25951 2534 25985 2568
rect 26023 2534 26032 2568
rect 26032 2534 26057 2568
rect 956 1674 960 1704
rect 960 1674 990 1704
rect 1028 1674 1062 1704
rect 1100 1699 25110 1703
rect 25149 1699 25183 1703
rect 25222 1699 25256 1703
rect 25295 1699 25329 1703
rect 25368 1699 25402 1703
rect 25441 1699 25475 1703
rect 25514 1699 25548 1703
rect 25587 1699 25621 1703
rect 25660 1699 25694 1703
rect 25733 1699 25767 1703
rect 25806 1699 25840 1703
rect 956 1670 990 1674
rect 1028 1670 1062 1674
rect 1100 1631 25110 1699
rect 25149 1669 25183 1699
rect 25222 1669 25256 1699
rect 25295 1669 25329 1699
rect 25368 1669 25402 1699
rect 25441 1669 25475 1699
rect 25514 1669 25548 1699
rect 25587 1669 25621 1699
rect 25660 1669 25694 1699
rect 25733 1669 25767 1699
rect 25806 1669 25814 1699
rect 25814 1669 25840 1699
rect 25879 1669 26032 2495
rect 956 1606 960 1631
rect 960 1606 990 1631
rect 956 1597 990 1606
rect 1028 1529 25182 1631
rect 25221 1597 25255 1631
rect 25294 1597 25328 1631
rect 25367 1597 25401 1631
rect 25440 1597 25474 1631
rect 25513 1597 25547 1631
rect 25586 1597 25620 1631
rect 25659 1597 25693 1631
rect 25732 1597 25766 1631
rect 25805 1597 25839 1631
rect 25878 1597 25882 1631
rect 25882 1597 25912 1631
rect 25951 1597 26032 1669
rect 26032 1597 26057 2495
rect 25221 1529 25255 1559
rect 25294 1529 25328 1559
rect 25367 1529 25401 1559
rect 25440 1529 25474 1559
rect 25513 1529 25547 1559
rect 25586 1529 25620 1559
rect 25659 1529 25693 1559
rect 25732 1529 25766 1559
rect 25805 1529 25839 1559
rect 25878 1529 25882 1559
rect 25882 1529 25912 1559
rect 1028 1525 25182 1529
rect 25221 1525 25255 1529
rect 25294 1525 25328 1529
rect 25367 1525 25401 1529
rect 25440 1525 25474 1529
rect 25513 1525 25547 1529
rect 25586 1525 25620 1529
rect 25659 1525 25693 1529
rect 25732 1525 25766 1529
rect 25805 1525 25839 1529
rect 25878 1525 25912 1529
rect 25951 1525 25985 1559
rect 26277 7705 26281 7739
rect 26281 7705 26311 7739
rect 26349 7703 26383 7737
rect 26421 7703 26451 7737
rect 26451 7703 26455 7737
rect 26277 7631 26281 7665
rect 26281 7631 26311 7665
rect 26349 7629 26383 7663
rect 26421 7629 26451 7663
rect 26451 7629 26455 7663
rect 26277 7557 26281 7591
rect 26281 7557 26311 7591
rect 26349 7556 26383 7590
rect 26421 7556 26451 7590
rect 26451 7556 26455 7590
rect 26277 7483 26281 7517
rect 26281 7483 26311 7517
rect 26349 7483 26383 7517
rect 26421 7483 26451 7517
rect 26451 7483 26455 7517
rect 26277 7373 26281 7407
rect 26281 7373 26311 7407
rect 26349 7373 26383 7407
rect 26421 7373 26451 7407
rect 26451 7373 26455 7407
rect 26277 7300 26281 7334
rect 26281 7300 26311 7334
rect 26349 7300 26383 7334
rect 26421 7300 26451 7334
rect 26451 7300 26455 7334
rect 26277 7227 26281 7261
rect 26281 7227 26311 7261
rect 26349 7227 26383 7261
rect 26421 7227 26451 7261
rect 26451 7227 26455 7261
rect 26277 7154 26281 7188
rect 26281 7154 26311 7188
rect 26349 7154 26383 7188
rect 26421 7154 26451 7188
rect 26451 7154 26455 7188
rect 26277 7081 26281 7115
rect 26281 7081 26311 7115
rect 26349 7081 26383 7115
rect 26421 7081 26451 7115
rect 26451 7081 26455 7115
rect 714 1475 744 1509
rect 744 1475 748 1509
rect 570 1403 574 1437
rect 574 1403 604 1437
rect 642 1403 676 1437
rect 714 1402 744 1436
rect 744 1402 748 1436
rect 570 1330 574 1364
rect 574 1330 604 1364
rect 642 1330 676 1364
rect 714 1329 744 1363
rect 744 1329 748 1363
rect 570 1257 574 1291
rect 574 1257 604 1291
rect 642 1257 676 1291
rect 714 1256 744 1290
rect 744 1256 748 1290
rect 570 1184 574 1218
rect 574 1184 604 1218
rect 642 1184 676 1218
rect 714 1183 744 1217
rect 744 1183 748 1217
rect 570 1111 574 1145
rect 574 1111 604 1145
rect 642 1111 676 1145
rect 714 1110 744 1144
rect 744 1110 748 1144
rect 570 1038 574 1072
rect 574 1038 604 1072
rect 642 1038 676 1072
rect 714 1037 744 1071
rect 744 1037 748 1071
rect 570 965 574 999
rect 574 965 604 999
rect 642 965 676 999
rect 714 964 744 998
rect 744 964 748 998
rect 570 892 574 926
rect 574 892 604 926
rect 642 892 676 926
rect 714 891 744 925
rect 744 891 748 925
rect 570 819 574 853
rect 574 819 604 853
rect 642 819 676 853
rect 714 818 744 852
rect 744 818 748 852
rect 570 746 574 780
rect 574 746 604 780
rect 642 746 676 780
rect 714 745 744 779
rect 744 745 748 779
rect 26277 2559 26281 7042
rect 26281 2559 26451 7042
rect 26277 2524 26349 2559
rect 26277 2490 26281 2524
rect 26281 2490 26315 2524
rect 26315 2491 26349 2524
rect 26349 2491 26451 2559
rect 26451 2491 26455 7042
rect 26315 2490 26455 2491
rect 26277 2456 26455 2490
rect 26277 2455 26349 2456
rect 26277 2421 26281 2455
rect 26281 2421 26315 2455
rect 26315 2422 26349 2455
rect 26349 2422 26383 2456
rect 26383 2422 26417 2456
rect 26417 2422 26451 2456
rect 26451 2422 26455 2456
rect 26315 2421 26455 2422
rect 26277 2387 26455 2421
rect 26277 2386 26349 2387
rect 26277 2352 26281 2386
rect 26281 2352 26315 2386
rect 26315 2353 26349 2386
rect 26349 2353 26383 2387
rect 26383 2353 26417 2387
rect 26417 2353 26451 2387
rect 26451 2353 26455 2387
rect 26315 2352 26455 2353
rect 26277 2318 26455 2352
rect 26277 2317 26349 2318
rect 26277 2283 26281 2317
rect 26281 2283 26315 2317
rect 26315 2284 26349 2317
rect 26349 2284 26383 2318
rect 26383 2284 26417 2318
rect 26417 2284 26451 2318
rect 26451 2284 26455 2318
rect 26315 2283 26455 2284
rect 26277 2249 26455 2283
rect 26277 2248 26349 2249
rect 26277 2214 26281 2248
rect 26281 2214 26315 2248
rect 26315 2215 26349 2248
rect 26349 2215 26383 2249
rect 26383 2215 26417 2249
rect 26417 2215 26451 2249
rect 26451 2215 26455 2249
rect 26315 2214 26455 2215
rect 26277 2180 26455 2214
rect 26277 2179 26349 2180
rect 26277 2145 26281 2179
rect 26281 2145 26315 2179
rect 26315 2146 26349 2179
rect 26349 2146 26383 2180
rect 26383 2146 26417 2180
rect 26417 2146 26451 2180
rect 26451 2146 26455 2180
rect 26315 2145 26455 2146
rect 26277 2111 26455 2145
rect 26277 2110 26349 2111
rect 26277 2076 26281 2110
rect 26281 2076 26315 2110
rect 26315 2077 26349 2110
rect 26349 2077 26383 2111
rect 26383 2077 26417 2111
rect 26417 2077 26451 2111
rect 26451 2077 26455 2111
rect 26315 2076 26455 2077
rect 26277 2042 26455 2076
rect 26277 2041 26349 2042
rect 26277 2007 26281 2041
rect 26281 2007 26315 2041
rect 26315 2008 26349 2041
rect 26349 2008 26383 2042
rect 26383 2008 26417 2042
rect 26417 2008 26451 2042
rect 26451 2008 26455 2042
rect 26315 2007 26455 2008
rect 26277 1973 26455 2007
rect 26277 1972 26349 1973
rect 26277 1938 26281 1972
rect 26281 1938 26315 1972
rect 26315 1939 26349 1972
rect 26349 1939 26383 1973
rect 26383 1939 26417 1973
rect 26417 1939 26451 1973
rect 26451 1939 26455 1973
rect 26315 1938 26455 1939
rect 26277 1904 26455 1938
rect 26277 1903 26349 1904
rect 26277 1869 26281 1903
rect 26281 1869 26315 1903
rect 26315 1870 26349 1903
rect 26349 1870 26383 1904
rect 26383 1870 26417 1904
rect 26417 1870 26451 1904
rect 26451 1870 26455 1904
rect 26315 1869 26455 1870
rect 26277 1835 26455 1869
rect 26277 1834 26349 1835
rect 26277 1800 26281 1834
rect 26281 1800 26315 1834
rect 26315 1801 26349 1834
rect 26349 1801 26383 1835
rect 26383 1801 26417 1835
rect 26417 1801 26451 1835
rect 26451 1801 26455 1835
rect 26315 1800 26455 1801
rect 26277 1766 26455 1800
rect 26277 1765 26349 1766
rect 26277 1731 26281 1765
rect 26281 1731 26315 1765
rect 26315 1732 26349 1765
rect 26349 1732 26383 1766
rect 26383 1732 26417 1766
rect 26417 1732 26451 1766
rect 26451 1732 26455 1766
rect 26315 1731 26455 1732
rect 26277 1697 26455 1731
rect 26277 1696 26349 1697
rect 26277 1662 26281 1696
rect 26281 1662 26315 1696
rect 26315 1663 26349 1696
rect 26349 1663 26383 1697
rect 26383 1663 26417 1697
rect 26417 1663 26451 1697
rect 26451 1663 26455 1697
rect 26315 1662 26455 1663
rect 26277 1628 26455 1662
rect 26277 1627 26349 1628
rect 26277 1593 26281 1627
rect 26281 1593 26315 1627
rect 26315 1594 26349 1627
rect 26349 1594 26383 1628
rect 26383 1594 26417 1628
rect 26417 1594 26451 1628
rect 26451 1594 26455 1628
rect 26315 1593 26455 1594
rect 26277 1559 26455 1593
rect 26277 1558 26349 1559
rect 26277 1524 26281 1558
rect 26281 1524 26315 1558
rect 26315 1525 26349 1558
rect 26349 1525 26383 1559
rect 26383 1525 26417 1559
rect 26417 1525 26451 1559
rect 26451 1525 26455 1559
rect 26315 1524 26455 1525
rect 26277 1490 26455 1524
rect 26277 1489 26349 1490
rect 26277 1455 26281 1489
rect 26281 1455 26315 1489
rect 26315 1456 26349 1489
rect 26349 1456 26383 1490
rect 26383 1456 26417 1490
rect 26417 1456 26451 1490
rect 26451 1456 26455 1490
rect 26315 1455 26455 1456
rect 26277 1421 26455 1455
rect 26277 1420 26349 1421
rect 26277 1386 26281 1420
rect 26281 1386 26315 1420
rect 26315 1387 26349 1420
rect 26349 1387 26383 1421
rect 26383 1387 26417 1421
rect 26417 1387 26451 1421
rect 26451 1387 26455 1421
rect 26315 1386 26455 1387
rect 26277 1352 26455 1386
rect 26277 1351 26349 1352
rect 26277 1317 26281 1351
rect 26281 1317 26315 1351
rect 26315 1318 26349 1351
rect 26349 1318 26383 1352
rect 26383 1318 26417 1352
rect 26417 1318 26451 1352
rect 26451 1318 26455 1352
rect 26315 1317 26455 1318
rect 26277 1283 26455 1317
rect 26277 1282 26349 1283
rect 26277 1248 26281 1282
rect 26281 1248 26315 1282
rect 26315 1249 26349 1282
rect 26349 1249 26383 1283
rect 26383 1249 26417 1283
rect 26417 1249 26451 1283
rect 26451 1249 26455 1283
rect 26315 1248 26455 1249
rect 26277 1214 26455 1248
rect 26277 1213 26349 1214
rect 26277 1179 26281 1213
rect 26281 1179 26315 1213
rect 26315 1180 26349 1213
rect 26349 1180 26383 1214
rect 26383 1180 26417 1214
rect 26417 1180 26451 1214
rect 26451 1180 26455 1214
rect 26315 1179 26455 1180
rect 26277 1145 26455 1179
rect 26277 1144 26349 1145
rect 26277 1110 26281 1144
rect 26281 1110 26315 1144
rect 26315 1111 26349 1144
rect 26349 1111 26383 1145
rect 26383 1111 26417 1145
rect 26417 1111 26451 1145
rect 26451 1111 26455 1145
rect 26315 1110 26455 1111
rect 26277 1076 26455 1110
rect 26277 1075 26349 1076
rect 26277 1041 26281 1075
rect 26281 1041 26315 1075
rect 26315 1042 26349 1075
rect 26349 1042 26383 1076
rect 26383 1042 26417 1076
rect 26417 1042 26451 1076
rect 26451 1042 26455 1076
rect 26315 1041 26455 1042
rect 26277 1007 26455 1041
rect 26277 1006 26349 1007
rect 26277 972 26281 1006
rect 26281 972 26315 1006
rect 26315 973 26349 1006
rect 26349 973 26383 1007
rect 26383 973 26417 1007
rect 26417 973 26451 1007
rect 26451 973 26455 1007
rect 26315 972 26455 973
rect 26277 938 26455 972
rect 26277 937 26349 938
rect 26277 903 26281 937
rect 26281 903 26315 937
rect 26315 904 26349 937
rect 26349 904 26383 938
rect 26383 904 26417 938
rect 26417 904 26451 938
rect 26451 904 26455 938
rect 26315 903 26455 904
rect 26277 869 26455 903
rect 26277 868 26349 869
rect 26277 834 26281 868
rect 26281 834 26315 868
rect 26315 835 26349 868
rect 26349 835 26383 869
rect 26383 835 26417 869
rect 26417 835 26451 869
rect 26451 835 26455 869
rect 26315 834 26455 835
rect 26277 800 26455 834
rect 26277 799 26349 800
rect 26277 765 26281 799
rect 26281 765 26315 799
rect 26315 766 26349 799
rect 26349 766 26383 800
rect 26383 766 26417 800
rect 26417 766 26451 800
rect 26451 766 26455 800
rect 26315 765 26455 766
rect 26277 731 26455 765
rect 26277 730 26349 731
rect 570 673 574 707
rect 574 673 604 707
rect 642 673 676 707
rect 714 696 744 706
rect 744 696 779 706
rect 779 696 813 706
rect 813 696 848 706
rect 848 696 882 706
rect 882 696 917 706
rect 714 662 917 696
rect 917 662 26092 706
rect 26131 672 26165 706
rect 26204 672 26238 706
rect 26277 672 26315 730
rect 26315 697 26349 730
rect 26349 697 26383 731
rect 26383 697 26417 731
rect 26417 697 26451 731
rect 26451 697 26455 731
rect 26315 672 26455 697
rect 26349 662 26455 672
rect 714 634 745 662
rect 570 628 574 634
rect 574 628 604 634
rect 642 628 676 634
rect 676 628 711 634
rect 711 628 745 634
rect 745 628 780 662
rect 780 628 814 662
rect 814 628 849 662
rect 849 634 26092 662
rect 570 600 604 628
rect 642 594 849 628
rect 642 560 676 594
rect 676 560 711 594
rect 711 560 745 594
rect 745 560 780 594
rect 780 560 814 594
rect 814 560 849 594
rect 849 560 26164 634
rect 26203 600 26237 634
rect 26276 600 26310 634
rect 26349 600 26383 662
rect 26383 628 26417 662
rect 26417 628 26451 662
rect 26451 628 26455 662
rect 26383 600 26455 628
rect 26203 560 26237 562
rect 26276 560 26310 562
rect 26349 560 26383 562
rect 642 528 26164 560
rect 26203 528 26237 560
rect 26276 528 26310 560
rect 26349 528 26383 560
rect 26680 8099 26684 8133
rect 26684 8099 26714 8133
rect 26752 8099 26786 8133
rect 26824 8099 26854 8133
rect 26854 8099 26858 8133
rect 26680 8020 26684 8054
rect 26684 8020 26714 8054
rect 26752 8020 26786 8054
rect 26824 8020 26854 8054
rect 26854 8020 26858 8054
rect 26680 7941 26684 7975
rect 26684 7941 26714 7975
rect 26752 7941 26786 7975
rect 26824 7941 26854 7975
rect 26854 7941 26858 7975
rect 26680 7862 26684 7896
rect 26684 7862 26714 7896
rect 26752 7862 26786 7896
rect 26824 7862 26854 7896
rect 26854 7862 26858 7896
rect 26680 7752 26684 7786
rect 26684 7752 26714 7786
rect 26752 7752 26786 7786
rect 26824 7752 26854 7786
rect 26854 7752 26858 7786
rect 26680 7679 26684 7713
rect 26684 7679 26714 7713
rect 26752 7679 26786 7713
rect 26824 7679 26854 7713
rect 26854 7679 26858 7713
rect 26680 7606 26684 7640
rect 26684 7606 26714 7640
rect 26752 7606 26786 7640
rect 26824 7606 26854 7640
rect 26854 7606 26858 7640
rect 26680 7533 26684 7567
rect 26684 7533 26714 7567
rect 26752 7533 26786 7567
rect 26824 7533 26854 7567
rect 26854 7533 26858 7567
rect 122 447 126 481
rect 126 447 156 481
rect 194 447 228 481
rect 266 446 296 480
rect 296 446 300 480
rect 122 374 126 408
rect 126 374 156 408
rect 194 374 228 408
rect 266 373 296 407
rect 296 373 300 407
rect 122 301 126 335
rect 126 301 156 335
rect 194 301 228 335
rect 266 262 296 334
rect 122 228 126 262
rect 126 228 156 262
rect 194 236 296 262
rect 296 236 22548 334
rect 22587 300 22621 334
rect 22660 300 22694 334
rect 22733 300 22767 334
rect 22806 300 22840 334
rect 22879 300 22913 334
rect 22952 300 22986 334
rect 23025 300 23059 334
rect 23098 300 23132 334
rect 23171 300 23205 334
rect 23244 300 23278 334
rect 23317 300 23351 334
rect 23390 300 23424 334
rect 23463 300 23497 334
rect 23536 300 23570 334
rect 23609 300 23643 334
rect 23682 300 23716 334
rect 23755 300 23789 334
rect 23828 300 23862 334
rect 23901 300 23935 334
rect 23974 300 24008 334
rect 24047 300 24081 334
rect 24120 300 24154 334
rect 24193 300 24227 334
rect 24266 300 24300 334
rect 24339 300 24373 334
rect 24412 300 24446 334
rect 24485 300 24519 334
rect 24558 300 24592 334
rect 24631 300 24665 334
rect 24704 300 24738 334
rect 24777 300 24811 334
rect 24850 300 24884 334
rect 24923 300 24957 334
rect 24996 300 25030 334
rect 25069 300 25103 334
rect 25142 300 25176 334
rect 25215 300 25249 334
rect 25288 300 25322 334
rect 25361 300 25395 334
rect 25434 300 25468 334
rect 25507 300 25541 334
rect 25580 300 25614 334
rect 25653 300 25687 334
rect 25726 300 25760 334
rect 25799 300 25833 334
rect 25872 300 25906 334
rect 25945 300 25979 334
rect 26018 300 26052 334
rect 26091 300 26125 334
rect 26164 300 26198 334
rect 26237 300 26271 334
rect 26310 300 26344 334
rect 26383 300 26417 334
rect 26456 300 26490 334
rect 26529 300 26563 334
rect 26602 300 26636 334
rect 22587 236 22621 262
rect 22660 236 22694 262
rect 22733 236 22767 262
rect 22806 236 22840 262
rect 22879 236 22913 262
rect 22952 236 22986 262
rect 23025 236 23059 262
rect 23098 236 23132 262
rect 23171 236 23205 262
rect 23244 236 23278 262
rect 23317 236 23351 262
rect 23390 236 23424 262
rect 23463 236 23497 262
rect 23536 236 23570 262
rect 23609 236 23643 262
rect 23682 236 23716 262
rect 23755 236 23789 262
rect 23828 236 23862 262
rect 23901 236 23935 262
rect 23974 236 24008 262
rect 24047 236 24081 262
rect 24120 236 24154 262
rect 24193 236 24227 262
rect 24266 236 24300 262
rect 24339 236 24373 262
rect 24412 236 24446 262
rect 24485 236 24519 262
rect 24558 236 24592 262
rect 24631 236 24665 262
rect 24704 236 24738 262
rect 24777 236 24811 262
rect 24850 236 24884 262
rect 24923 236 24957 262
rect 24996 236 25030 262
rect 25069 236 25103 262
rect 25142 236 25176 262
rect 25215 236 25249 262
rect 25288 236 25322 262
rect 25361 236 25395 262
rect 25434 236 25468 262
rect 25507 236 25541 262
rect 25580 236 25614 262
rect 25653 236 25687 262
rect 25726 236 25760 262
rect 25799 236 25833 262
rect 25872 236 25906 262
rect 25945 236 25979 262
rect 26018 236 26052 262
rect 26091 236 26125 262
rect 26164 236 26198 262
rect 26237 236 26271 262
rect 26310 236 26344 262
rect 26383 236 26417 262
rect 26456 236 26490 262
rect 26529 236 26563 262
rect 26602 236 26636 262
rect 26680 236 26684 7494
rect 26684 236 26854 7494
rect 194 156 364 236
rect 364 202 399 236
rect 399 202 433 236
rect 433 202 468 236
rect 468 202 502 236
rect 502 202 537 236
rect 537 202 571 236
rect 571 202 606 236
rect 606 202 640 236
rect 640 202 675 236
rect 675 202 709 236
rect 709 202 744 236
rect 744 202 778 236
rect 778 202 813 236
rect 813 202 847 236
rect 847 202 882 236
rect 882 202 916 236
rect 916 202 951 236
rect 951 202 985 236
rect 985 202 1020 236
rect 1020 202 1054 236
rect 1054 202 1089 236
rect 1089 202 1123 236
rect 1123 202 1158 236
rect 1158 202 1192 236
rect 1192 202 1227 236
rect 1227 202 1261 236
rect 1261 202 1296 236
rect 1296 202 1330 236
rect 1330 202 1365 236
rect 1365 202 1399 236
rect 1399 202 1434 236
rect 1434 202 1468 236
rect 1468 202 1503 236
rect 1503 202 1537 236
rect 1537 202 1572 236
rect 1572 202 1606 236
rect 1606 202 1641 236
rect 1641 202 1675 236
rect 1675 202 1710 236
rect 1710 202 1744 236
rect 1744 202 1779 236
rect 1779 202 1813 236
rect 1813 202 1848 236
rect 1848 202 1882 236
rect 1882 202 1917 236
rect 1917 202 1951 236
rect 1951 202 1986 236
rect 1986 202 2020 236
rect 2020 202 2055 236
rect 2055 202 2089 236
rect 2089 202 2124 236
rect 2124 202 2158 236
rect 2158 202 2193 236
rect 2193 202 2227 236
rect 2227 202 2262 236
rect 2262 202 2296 236
rect 2296 202 2331 236
rect 2331 202 2365 236
rect 2365 202 2400 236
rect 2400 202 2434 236
rect 2434 202 2469 236
rect 2469 202 2503 236
rect 2503 202 2538 236
rect 2538 202 2572 236
rect 2572 202 2607 236
rect 2607 202 2641 236
rect 2641 202 2676 236
rect 2676 202 2710 236
rect 2710 202 2745 236
rect 2745 202 2779 236
rect 2779 202 2814 236
rect 2814 202 2848 236
rect 2848 202 2883 236
rect 2883 202 2917 236
rect 2917 202 2952 236
rect 364 168 2952 202
rect 364 156 399 168
rect 399 156 433 168
rect 433 156 468 168
rect 468 156 502 168
rect 502 156 537 168
rect 537 156 571 168
rect 571 156 606 168
rect 606 156 640 168
rect 640 156 675 168
rect 675 156 709 168
rect 709 156 744 168
rect 744 156 778 168
rect 778 156 813 168
rect 813 156 847 168
rect 847 156 882 168
rect 882 156 916 168
rect 916 156 951 168
rect 951 156 985 168
rect 985 156 1020 168
rect 1020 156 1054 168
rect 1054 156 1089 168
rect 1089 156 1123 168
rect 1123 156 1158 168
rect 1158 156 1192 168
rect 1192 156 1227 168
rect 1227 156 1261 168
rect 1261 156 1296 168
rect 1296 156 1330 168
rect 1330 156 1365 168
rect 1365 156 1399 168
rect 1399 156 1434 168
rect 1434 156 1468 168
rect 1468 156 1503 168
rect 1503 156 1537 168
rect 1537 156 1572 168
rect 1572 156 1606 168
rect 1606 156 1641 168
rect 1641 156 1675 168
rect 1675 156 1710 168
rect 1710 156 1744 168
rect 1744 156 1779 168
rect 1779 156 1813 168
rect 1813 156 1848 168
rect 1848 156 1882 168
rect 1882 156 1917 168
rect 1917 156 1951 168
rect 1951 156 1986 168
rect 1986 156 2020 168
rect 2020 156 2055 168
rect 2055 156 2089 168
rect 2089 156 2124 168
rect 2124 156 2158 168
rect 2158 156 2193 168
rect 2193 156 2227 168
rect 2227 156 2262 168
rect 2262 156 2296 168
rect 2296 156 2331 168
rect 2331 156 2365 168
rect 2365 156 2400 168
rect 2400 156 2434 168
rect 2434 156 2469 168
rect 2469 156 2503 168
rect 2503 156 2538 168
rect 2538 156 2572 168
rect 2572 156 2607 168
rect 2607 156 2641 168
rect 2641 156 2676 168
rect 2676 156 2710 168
rect 2710 156 2745 168
rect 2745 156 2779 168
rect 2779 156 2814 168
rect 2814 156 2848 168
rect 2848 156 2883 168
rect 2883 156 2917 168
rect 2917 156 2952 168
rect 2952 156 22548 236
rect 22587 228 22621 236
rect 22660 228 22694 236
rect 22733 228 22767 236
rect 22806 228 22840 236
rect 22879 228 22913 236
rect 22952 228 22986 236
rect 23025 228 23059 236
rect 23098 228 23132 236
rect 23171 228 23205 236
rect 23244 228 23278 236
rect 23317 228 23351 236
rect 23390 228 23424 236
rect 23463 228 23497 236
rect 23536 228 23570 236
rect 23609 228 23643 236
rect 23682 228 23716 236
rect 23755 228 23789 236
rect 23828 228 23862 236
rect 23901 228 23935 236
rect 23974 228 24008 236
rect 24047 228 24081 236
rect 24120 228 24154 236
rect 24193 228 24227 236
rect 24266 228 24300 236
rect 24339 228 24373 236
rect 24412 228 24446 236
rect 24485 228 24519 236
rect 24558 228 24592 236
rect 24631 228 24665 236
rect 24704 228 24738 236
rect 24777 228 24811 236
rect 24850 228 24884 236
rect 24923 228 24957 236
rect 24996 228 25030 236
rect 25069 228 25103 236
rect 25142 228 25176 236
rect 25215 228 25249 236
rect 25288 228 25322 236
rect 25361 228 25395 236
rect 25434 228 25468 236
rect 25507 228 25541 236
rect 25580 228 25614 236
rect 25653 228 25687 236
rect 25726 228 25760 236
rect 25799 228 25833 236
rect 25872 228 25906 236
rect 25945 228 25979 236
rect 26018 228 26052 236
rect 26091 228 26125 236
rect 26164 228 26198 236
rect 26237 228 26271 236
rect 26310 228 26344 236
rect 26383 228 26417 236
rect 26456 228 26490 236
rect 26529 228 26563 236
rect 26602 228 26636 236
rect 22587 156 22621 190
rect 22660 156 22694 190
rect 22733 156 22767 190
rect 22806 156 22840 190
rect 22879 156 22913 190
rect 22952 156 22986 190
rect 23025 156 23059 190
rect 23098 156 23132 190
rect 23171 156 23205 190
rect 23244 156 23278 190
rect 23317 156 23351 190
rect 23390 156 23424 190
rect 23463 156 23497 190
rect 23536 156 23570 190
rect 23609 156 23643 190
rect 23682 156 23716 190
rect 23755 156 23789 190
rect 23828 156 23862 190
rect 23901 156 23935 190
rect 23974 156 24008 190
rect 24047 156 24081 190
rect 24120 156 24154 190
rect 24193 156 24227 190
rect 24266 156 24300 190
rect 24339 156 24373 190
rect 24412 156 24446 190
rect 24485 156 24519 190
rect 24558 156 24592 190
rect 24631 156 24665 190
rect 24704 156 24738 190
rect 24777 156 24811 190
rect 24850 156 24884 190
rect 24923 156 24957 190
rect 24996 156 25030 190
rect 25069 156 25103 190
rect 25142 156 25176 190
rect 25215 156 25249 190
rect 25288 156 25322 190
rect 25361 156 25395 190
rect 25434 156 25468 190
rect 25507 156 25541 190
rect 25580 156 25614 190
rect 25653 156 25687 190
rect 25726 156 25760 190
rect 25799 156 25833 190
rect 25872 156 25906 190
rect 25945 156 25979 190
rect 26018 156 26052 190
rect 26091 156 26125 190
rect 26164 156 26198 190
rect 26237 156 26271 190
rect 26310 156 26344 190
rect 26383 156 26417 190
rect 26456 156 26490 190
rect 26529 156 26563 190
rect 26602 156 26636 190
rect 26680 188 26854 236
rect 26854 188 26858 7494
<< metal1 >>
rect 116 8484 26864 8490
rect 116 8450 194 8484
rect 228 8450 267 8484
rect 301 8450 340 8484
rect 374 8450 413 8484
rect 447 8450 486 8484
rect 520 8450 559 8484
rect 593 8450 632 8484
rect 666 8450 705 8484
rect 739 8450 778 8484
rect 812 8450 851 8484
rect 885 8450 924 8484
rect 958 8450 997 8484
rect 1031 8450 1070 8484
rect 1104 8450 1143 8484
rect 1177 8450 1216 8484
rect 1250 8450 1289 8484
rect 1323 8450 1362 8484
rect 1396 8450 1435 8484
rect 1469 8450 1508 8484
rect 1542 8450 1581 8484
rect 1615 8450 1654 8484
rect 1688 8450 1727 8484
rect 1761 8450 1800 8484
rect 1834 8450 1873 8484
rect 1907 8450 1946 8484
rect 1980 8450 2019 8484
rect 2053 8450 2092 8484
rect 2126 8450 2165 8484
rect 2199 8450 2238 8484
rect 2272 8450 2311 8484
rect 2345 8450 2384 8484
rect 2418 8450 2457 8484
rect 2491 8450 2530 8484
rect 2564 8450 2603 8484
rect 2637 8450 2676 8484
rect 2710 8450 2749 8484
rect 2783 8450 2822 8484
rect 2856 8450 2895 8484
rect 2929 8450 2968 8484
rect 3002 8450 3041 8484
rect 3075 8450 3114 8484
rect 3148 8450 3187 8484
rect 3221 8450 3260 8484
rect 3294 8450 3333 8484
rect 3367 8450 3406 8484
rect 3440 8450 3479 8484
rect 3513 8450 3552 8484
rect 3586 8450 3625 8484
rect 3659 8450 3698 8484
rect 3732 8450 3771 8484
rect 3805 8450 3844 8484
rect 3878 8450 3917 8484
rect 3951 8450 3990 8484
rect 4024 8450 4063 8484
rect 4097 8450 4136 8484
rect 4170 8450 4209 8484
rect 4243 8450 4282 8484
rect 116 8412 4282 8450
rect 116 1250 122 8412
rect 228 8378 267 8412
rect 301 8378 340 8412
rect 374 8378 413 8412
rect 447 8378 486 8412
rect 520 8378 559 8412
rect 593 8378 632 8412
rect 666 8378 705 8412
rect 739 8378 778 8412
rect 812 8378 851 8412
rect 885 8378 924 8412
rect 958 8378 997 8412
rect 1031 8378 1070 8412
rect 1104 8378 1143 8412
rect 1177 8378 1216 8412
rect 1250 8378 1289 8412
rect 1323 8378 1362 8412
rect 1396 8378 1435 8412
rect 1469 8378 1508 8412
rect 1542 8378 1581 8412
rect 1615 8378 1654 8412
rect 1688 8378 1727 8412
rect 1761 8378 1800 8412
rect 1834 8378 1873 8412
rect 1907 8378 1946 8412
rect 1980 8378 2019 8412
rect 2053 8378 2092 8412
rect 2126 8378 2165 8412
rect 2199 8378 2238 8412
rect 2272 8378 2311 8412
rect 2345 8378 2384 8412
rect 2418 8378 2457 8412
rect 2491 8378 2530 8412
rect 2564 8378 2603 8412
rect 2637 8378 2676 8412
rect 2710 8378 2749 8412
rect 2783 8378 2822 8412
rect 2856 8378 2895 8412
rect 2929 8378 2968 8412
rect 3002 8378 3041 8412
rect 3075 8378 3114 8412
rect 3148 8378 3187 8412
rect 3221 8378 3260 8412
rect 3294 8378 3333 8412
rect 3367 8378 3406 8412
rect 3440 8378 3479 8412
rect 3513 8378 3552 8412
rect 3586 8378 3625 8412
rect 3659 8378 3698 8412
rect 3732 8378 3771 8412
rect 3805 8378 3844 8412
rect 3878 8378 3917 8412
rect 3951 8378 3990 8412
rect 4024 8378 4063 8412
rect 4097 8378 4136 8412
rect 4170 8378 4209 8412
rect 4243 8378 4282 8412
rect 26636 8452 26864 8484
rect 26636 8418 26680 8452
rect 26714 8418 26752 8452
rect 26786 8418 26824 8452
rect 26858 8418 26864 8452
rect 228 8340 4354 8378
rect 300 8306 339 8340
rect 373 8306 412 8340
rect 446 8306 485 8340
rect 519 8306 558 8340
rect 592 8306 631 8340
rect 665 8306 704 8340
rect 738 8306 777 8340
rect 811 8306 850 8340
rect 884 8306 923 8340
rect 957 8306 996 8340
rect 1030 8306 1069 8340
rect 1103 8306 1142 8340
rect 1176 8306 1215 8340
rect 1249 8306 1288 8340
rect 1322 8306 1361 8340
rect 1395 8306 1434 8340
rect 1468 8306 1507 8340
rect 1541 8306 1580 8340
rect 1614 8306 1653 8340
rect 1687 8306 1726 8340
rect 1760 8306 1799 8340
rect 1833 8306 1872 8340
rect 1906 8306 1945 8340
rect 1979 8306 2018 8340
rect 2052 8306 2091 8340
rect 2125 8306 2164 8340
rect 2198 8306 2237 8340
rect 2271 8306 2310 8340
rect 2344 8306 2383 8340
rect 2417 8306 2456 8340
rect 2490 8306 2529 8340
rect 2563 8306 2602 8340
rect 2636 8306 2675 8340
rect 2709 8306 2748 8340
rect 2782 8306 2821 8340
rect 2855 8306 2894 8340
rect 2928 8306 2967 8340
rect 3001 8306 3040 8340
rect 3074 8306 3113 8340
rect 3147 8306 3186 8340
rect 3220 8306 3259 8340
rect 3293 8306 3332 8340
rect 3366 8306 3405 8340
rect 3439 8306 3478 8340
rect 3512 8306 3551 8340
rect 3585 8306 3624 8340
rect 3658 8306 3697 8340
rect 3731 8306 3770 8340
rect 3804 8306 3843 8340
rect 3877 8306 3916 8340
rect 3950 8306 3989 8340
rect 4023 8306 4062 8340
rect 4096 8306 4135 8340
rect 4169 8306 4208 8340
rect 4242 8306 4281 8340
rect 4315 8306 4354 8340
rect 26636 8372 26864 8418
rect 26636 8338 26680 8372
rect 26714 8338 26752 8372
rect 26786 8338 26824 8372
rect 26858 8338 26864 8372
rect 26636 8306 26864 8338
rect 300 8300 26864 8306
rect 300 8292 356 8300
tri 356 8292 364 8300 nw
tri 26616 8292 26624 8300 ne
rect 26624 8292 26864 8300
rect 300 8258 322 8292
tri 322 8258 356 8292 nw
tri 26624 8258 26658 8292 ne
rect 26658 8258 26680 8292
rect 26714 8258 26752 8292
rect 26786 8258 26824 8292
rect 26858 8258 26864 8292
rect 300 1322 306 8258
tri 306 8242 322 8258 nw
tri 26658 8242 26674 8258 ne
rect 26674 8212 26864 8258
rect 26674 8178 26680 8212
rect 26714 8178 26752 8212
rect 26786 8178 26824 8212
rect 26858 8178 26864 8212
rect 26674 8133 26864 8178
rect 228 1283 306 1322
rect 228 1250 266 1283
rect 116 1249 266 1250
rect 300 1249 306 1283
rect 116 1211 306 1249
rect 116 1177 122 1211
rect 156 1177 194 1211
rect 228 1210 306 1211
rect 228 1177 266 1210
rect 116 1176 266 1177
rect 300 1176 306 1210
rect 116 1138 306 1176
rect 116 1104 122 1138
rect 156 1104 194 1138
rect 228 1137 306 1138
rect 228 1104 266 1137
rect 116 1103 266 1104
rect 300 1103 306 1137
rect 116 1065 306 1103
rect 116 1031 122 1065
rect 156 1031 194 1065
rect 228 1064 306 1065
rect 228 1031 266 1064
rect 116 1030 266 1031
rect 300 1030 306 1064
rect 116 992 306 1030
rect 116 958 122 992
rect 156 958 194 992
rect 228 991 306 992
rect 228 958 266 991
rect 116 957 266 958
rect 300 957 306 991
rect 116 919 306 957
rect 116 885 122 919
rect 156 885 194 919
rect 228 918 306 919
rect 228 885 266 918
rect 116 884 266 885
rect 300 884 306 918
rect 116 846 306 884
rect 116 812 122 846
rect 156 812 194 846
rect 228 845 306 846
rect 228 812 266 845
rect 116 811 266 812
rect 300 811 306 845
rect 116 773 306 811
rect 116 739 122 773
rect 156 739 194 773
rect 228 772 306 773
rect 228 739 266 772
rect 116 738 266 739
rect 300 738 306 772
rect 116 700 306 738
rect 116 666 122 700
rect 156 666 194 700
rect 228 699 306 700
rect 228 666 266 699
rect 116 665 266 666
rect 300 665 306 699
rect 116 627 306 665
rect 116 593 122 627
rect 156 593 194 627
rect 228 626 306 627
rect 228 593 266 626
rect 116 592 266 593
rect 300 592 306 626
rect 116 554 306 592
rect 116 520 122 554
rect 156 520 194 554
rect 228 553 306 554
rect 228 520 266 553
rect 116 519 266 520
rect 300 519 306 553
rect 564 8105 26461 8111
rect 564 8071 642 8105
rect 676 8071 715 8105
rect 749 8071 788 8105
rect 822 8071 861 8105
rect 564 8033 861 8071
rect 564 4615 570 8033
rect 676 7999 715 8033
rect 749 7999 788 8033
rect 822 7999 861 8033
rect 26383 8033 26461 8105
rect 26383 7999 26421 8033
rect 26455 7999 26461 8033
rect 676 7961 933 7999
rect 748 7927 787 7961
rect 821 7927 860 7961
rect 894 7927 933 7961
rect 26311 7959 26461 7999
rect 26311 7927 26349 7959
rect 748 7925 26349 7927
rect 26383 7925 26421 7959
rect 26455 7925 26461 7959
rect 748 7921 26461 7925
rect 748 7896 795 7921
tri 795 7896 820 7921 nw
tri 26205 7896 26230 7921 ne
rect 26230 7896 26461 7921
rect 748 7887 786 7896
tri 786 7887 795 7896 nw
tri 26230 7887 26239 7896 ne
rect 26239 7887 26461 7896
rect 748 4687 754 7887
tri 754 7855 786 7887 nw
tri 26239 7855 26271 7887 ne
rect 26271 7853 26277 7887
rect 26311 7885 26461 7887
rect 26311 7853 26349 7885
rect 26271 7851 26349 7853
rect 26383 7851 26421 7885
rect 26455 7851 26461 7885
rect 26271 7813 26461 7851
rect 26271 7779 26277 7813
rect 26311 7811 26461 7813
rect 26311 7779 26349 7811
rect 26271 7777 26349 7779
rect 26383 7777 26421 7811
rect 26455 7777 26461 7811
rect 26271 7739 26461 7777
rect 676 4648 754 4687
rect 676 4615 714 4648
rect 564 4614 714 4615
rect 748 4614 754 4648
rect 564 4576 754 4614
rect 564 4542 570 4576
rect 604 4542 642 4576
rect 676 4575 754 4576
rect 676 4542 714 4575
rect 564 4541 714 4542
rect 748 4541 754 4575
rect 564 4503 754 4541
rect 564 4469 570 4503
rect 604 4469 642 4503
rect 676 4502 754 4503
rect 676 4469 714 4502
rect 564 4468 714 4469
rect 748 4468 754 4502
rect 564 4430 754 4468
rect 564 4396 570 4430
rect 604 4396 642 4430
rect 676 4429 754 4430
rect 676 4396 714 4429
rect 564 4395 714 4396
rect 748 4395 754 4429
rect 564 4357 754 4395
rect 564 4323 570 4357
rect 604 4323 642 4357
rect 676 4356 754 4357
rect 676 4323 714 4356
rect 564 4322 714 4323
rect 748 4322 754 4356
rect 564 4284 754 4322
rect 564 4250 570 4284
rect 604 4250 642 4284
rect 676 4283 754 4284
rect 676 4250 714 4283
rect 564 4249 714 4250
rect 748 4249 754 4283
rect 564 4211 754 4249
rect 564 4177 570 4211
rect 604 4177 642 4211
rect 676 4210 754 4211
rect 676 4177 714 4210
rect 564 4176 714 4177
rect 748 4176 754 4210
rect 564 4138 754 4176
rect 564 4104 570 4138
rect 604 4104 642 4138
rect 676 4137 754 4138
rect 676 4104 714 4137
rect 564 4103 714 4104
rect 748 4103 754 4137
rect 564 4065 754 4103
rect 564 4031 570 4065
rect 604 4031 642 4065
rect 676 4064 754 4065
rect 676 4031 714 4064
rect 564 4030 714 4031
rect 748 4030 754 4064
rect 564 3992 754 4030
rect 564 3958 570 3992
rect 604 3958 642 3992
rect 676 3991 754 3992
rect 676 3958 714 3991
rect 564 3957 714 3958
rect 748 3957 754 3991
rect 564 3919 754 3957
rect 564 3885 570 3919
rect 604 3885 642 3919
rect 676 3918 754 3919
rect 676 3885 714 3918
rect 564 3884 714 3885
rect 748 3884 754 3918
rect 564 3846 754 3884
rect 564 3812 570 3846
rect 604 3812 642 3846
rect 676 3845 754 3846
rect 676 3812 714 3845
rect 564 3811 714 3812
rect 748 3811 754 3845
rect 564 3773 754 3811
rect 564 3739 570 3773
rect 604 3739 642 3773
rect 676 3772 754 3773
rect 676 3739 714 3772
rect 564 3738 714 3739
rect 748 3738 754 3772
rect 564 3700 754 3738
rect 564 3666 570 3700
rect 604 3666 642 3700
rect 676 3699 754 3700
rect 676 3666 714 3699
rect 564 3665 714 3666
rect 748 3665 754 3699
rect 564 3627 754 3665
rect 564 3593 570 3627
rect 604 3593 642 3627
rect 676 3626 754 3627
rect 676 3593 714 3626
rect 564 3592 714 3593
rect 748 3592 754 3626
rect 564 3554 754 3592
rect 564 3520 570 3554
rect 604 3520 642 3554
rect 676 3553 754 3554
rect 676 3520 714 3553
rect 564 3519 714 3520
rect 748 3519 754 3553
rect 564 3481 754 3519
rect 564 3447 570 3481
rect 604 3447 642 3481
rect 676 3480 754 3481
rect 676 3447 714 3480
rect 564 3446 714 3447
rect 748 3446 754 3480
rect 564 3408 754 3446
rect 564 3374 570 3408
rect 604 3374 642 3408
rect 676 3407 754 3408
rect 676 3374 714 3407
rect 564 3373 714 3374
rect 748 3373 754 3407
rect 564 3335 754 3373
rect 564 3301 570 3335
rect 604 3301 642 3335
rect 676 3334 754 3335
rect 676 3301 714 3334
rect 564 3300 714 3301
rect 748 3300 754 3334
rect 564 3262 754 3300
rect 564 3228 570 3262
rect 604 3228 642 3262
rect 676 3261 754 3262
rect 676 3228 714 3261
rect 564 3227 714 3228
rect 748 3227 754 3261
rect 564 3189 754 3227
rect 564 3155 570 3189
rect 604 3155 642 3189
rect 676 3188 754 3189
rect 676 3155 714 3188
rect 564 3154 714 3155
rect 748 3154 754 3188
rect 564 3116 754 3154
rect 564 3082 570 3116
rect 604 3082 642 3116
rect 676 3115 754 3116
rect 676 3082 714 3115
rect 564 3081 714 3082
rect 748 3081 754 3115
rect 564 3043 754 3081
rect 564 3009 570 3043
rect 604 3009 642 3043
rect 676 3042 754 3043
rect 676 3009 714 3042
rect 564 3008 714 3009
rect 748 3008 754 3042
rect 564 2970 754 3008
rect 564 2936 570 2970
rect 604 2936 642 2970
rect 676 2969 754 2970
rect 676 2936 714 2969
rect 564 2935 714 2936
rect 748 2935 754 2969
rect 564 2897 754 2935
rect 564 2863 570 2897
rect 604 2863 642 2897
rect 676 2896 754 2897
rect 676 2863 714 2896
rect 564 2862 714 2863
rect 748 2862 754 2896
rect 564 2824 754 2862
rect 564 2790 570 2824
rect 604 2790 642 2824
rect 676 2823 754 2824
rect 676 2790 714 2823
rect 564 2789 714 2790
rect 748 2789 754 2823
rect 564 2751 754 2789
rect 564 2717 570 2751
rect 604 2717 642 2751
rect 676 2750 754 2751
rect 676 2717 714 2750
rect 564 2716 714 2717
rect 748 2716 754 2750
rect 564 2678 754 2716
rect 564 2644 570 2678
rect 604 2644 642 2678
rect 676 2677 754 2678
rect 676 2644 714 2677
rect 564 2643 714 2644
rect 748 2643 754 2677
rect 564 2605 754 2643
rect 564 2571 570 2605
rect 604 2571 642 2605
rect 676 2604 754 2605
rect 676 2571 714 2604
rect 564 2570 714 2571
rect 748 2570 754 2604
rect 564 2532 754 2570
rect 564 2498 570 2532
rect 604 2498 642 2532
rect 676 2531 754 2532
rect 676 2498 714 2531
rect 564 2497 714 2498
rect 748 2497 754 2531
rect 564 2459 754 2497
rect 564 2425 570 2459
rect 604 2425 642 2459
rect 676 2458 754 2459
rect 676 2425 714 2458
rect 564 2424 714 2425
rect 748 2424 754 2458
rect 564 2386 754 2424
rect 564 2352 570 2386
rect 604 2352 642 2386
rect 676 2385 754 2386
rect 676 2352 714 2385
rect 564 2351 714 2352
rect 748 2351 754 2385
rect 564 2313 754 2351
rect 564 2279 570 2313
rect 604 2279 642 2313
rect 676 2312 754 2313
rect 676 2279 714 2312
rect 564 2278 714 2279
rect 748 2278 754 2312
rect 564 2240 754 2278
rect 564 2206 570 2240
rect 604 2206 642 2240
rect 676 2239 754 2240
rect 676 2206 714 2239
rect 564 2205 714 2206
rect 748 2205 754 2239
rect 564 2167 754 2205
rect 564 2133 570 2167
rect 604 2133 642 2167
rect 676 2166 754 2167
rect 676 2133 714 2166
rect 564 2132 714 2133
rect 748 2132 754 2166
rect 564 2094 754 2132
rect 564 2060 570 2094
rect 604 2060 642 2094
rect 676 2093 754 2094
rect 676 2060 714 2093
rect 564 2059 714 2060
rect 748 2059 754 2093
rect 564 2021 754 2059
rect 564 1987 570 2021
rect 604 1987 642 2021
rect 676 2020 754 2021
rect 676 1987 714 2020
rect 564 1986 714 1987
rect 748 1986 754 2020
rect 564 1948 754 1986
rect 564 1914 570 1948
rect 604 1914 642 1948
rect 676 1947 754 1948
rect 676 1914 714 1947
rect 564 1913 714 1914
rect 748 1913 754 1947
rect 564 1875 754 1913
rect 564 1841 570 1875
rect 604 1841 642 1875
rect 676 1874 754 1875
rect 676 1841 714 1874
rect 564 1840 714 1841
rect 748 1840 754 1874
rect 564 1802 754 1840
rect 564 1768 570 1802
rect 604 1768 642 1802
rect 676 1801 754 1802
rect 676 1768 714 1801
rect 564 1767 714 1768
rect 748 1767 754 1801
rect 564 1729 754 1767
rect 564 1695 570 1729
rect 604 1695 642 1729
rect 676 1728 754 1729
rect 676 1695 714 1728
rect 564 1694 714 1695
rect 748 1694 754 1728
rect 564 1656 754 1694
rect 564 1622 570 1656
rect 604 1622 642 1656
rect 676 1655 754 1656
rect 676 1622 714 1655
rect 564 1621 714 1622
rect 748 1621 754 1655
rect 564 1583 754 1621
rect 564 1549 570 1583
rect 604 1549 642 1583
rect 676 1582 754 1583
rect 676 1549 714 1582
rect 564 1548 714 1549
rect 748 1548 754 1582
rect 564 1510 754 1548
rect 950 7719 26063 7725
rect 950 7685 1028 7719
rect 1062 7685 1101 7719
rect 1135 7685 1174 7719
rect 1208 7685 1247 7719
rect 1281 7685 1320 7719
rect 1354 7685 1393 7719
rect 1427 7685 1466 7719
rect 1500 7685 1539 7719
rect 1573 7685 1612 7719
rect 1646 7685 1685 7719
rect 1719 7685 1758 7719
rect 1792 7685 1831 7719
rect 950 7647 1831 7685
rect 950 4517 956 7647
rect 1062 7613 1101 7647
rect 1135 7613 1174 7647
rect 1208 7613 1247 7647
rect 1281 7613 1320 7647
rect 1354 7613 1393 7647
rect 1427 7613 1466 7647
rect 1500 7613 1539 7647
rect 1573 7613 1612 7647
rect 1646 7613 1685 7647
rect 1719 7613 1758 7647
rect 1792 7613 1831 7647
rect 25985 7647 26063 7719
rect 25985 7613 26023 7647
rect 26057 7613 26063 7647
rect 1062 7575 1903 7613
rect 1134 7541 1173 7575
rect 1207 7541 1246 7575
rect 1280 7541 1319 7575
rect 1353 7541 1392 7575
rect 1426 7541 1465 7575
rect 1499 7541 1538 7575
rect 1572 7541 1611 7575
rect 1645 7541 1684 7575
rect 1718 7541 1757 7575
rect 1791 7541 1830 7575
rect 1864 7541 1903 7575
rect 25913 7573 26063 7613
rect 25913 7541 25951 7573
rect 1134 7539 25951 7541
rect 25985 7539 26023 7573
rect 26057 7539 26063 7573
rect 1134 7535 26063 7539
rect 1134 7533 1172 7535
tri 1172 7533 1174 7535 nw
tri 25821 7533 25823 7535 ne
rect 25823 7533 26063 7535
rect 1134 7517 1156 7533
tri 1156 7517 1172 7533 nw
tri 25823 7517 25839 7533 ne
rect 25839 7517 26063 7533
rect 1134 4589 1140 7517
tri 1140 7501 1156 7517 nw
tri 25839 7501 25855 7517 ne
rect 25855 7501 26063 7517
tri 25855 7483 25873 7501 ne
rect 25873 7467 25879 7501
rect 25913 7499 26063 7501
rect 25913 7467 25951 7499
rect 25873 7465 25951 7467
rect 25985 7465 26023 7499
rect 26057 7465 26063 7499
rect 25873 7427 26063 7465
rect 1284 7393 1305 7416
tri 1305 7393 1328 7416 nw
rect 25873 7393 25879 7427
rect 25913 7425 26063 7427
rect 25913 7393 25951 7425
rect 1284 7391 1303 7393
tri 1303 7391 1305 7393 nw
rect 25873 7391 25951 7393
rect 25985 7391 26023 7425
rect 26057 7391 26063 7425
rect 1284 7373 1285 7391
tri 1285 7373 1303 7391 nw
tri 1284 7372 1285 7373 nw
rect 1062 4550 1140 4589
rect 1062 4517 1100 4550
rect 950 4516 1100 4517
rect 1134 4516 1140 4550
rect 950 4478 1140 4516
rect 950 4444 956 4478
rect 990 4444 1028 4478
rect 1062 4477 1140 4478
rect 1062 4444 1100 4477
rect 950 4443 1100 4444
rect 1134 4443 1140 4477
rect 950 4405 1140 4443
rect 950 4371 956 4405
rect 990 4371 1028 4405
rect 1062 4404 1140 4405
rect 1062 4371 1100 4404
rect 950 4370 1100 4371
rect 1134 4370 1140 4404
rect 950 4332 1140 4370
rect 950 4298 956 4332
rect 990 4298 1028 4332
rect 1062 4331 1140 4332
rect 1062 4298 1100 4331
rect 950 4297 1100 4298
rect 1134 4297 1140 4331
rect 950 4259 1140 4297
rect 950 4225 956 4259
rect 990 4225 1028 4259
rect 1062 4258 1140 4259
rect 1062 4225 1100 4258
rect 950 4224 1100 4225
rect 1134 4224 1140 4258
rect 950 4186 1140 4224
rect 950 4152 956 4186
rect 990 4152 1028 4186
rect 1062 4185 1140 4186
rect 1062 4152 1100 4185
rect 950 4151 1100 4152
rect 1134 4151 1140 4185
rect 950 4113 1140 4151
rect 950 4079 956 4113
rect 990 4079 1028 4113
rect 1062 4112 1140 4113
rect 1062 4079 1100 4112
rect 950 4078 1100 4079
rect 1134 4078 1140 4112
rect 950 4040 1140 4078
rect 950 4006 956 4040
rect 990 4006 1028 4040
rect 1062 4039 1140 4040
rect 1062 4006 1100 4039
rect 950 4005 1100 4006
rect 1134 4005 1140 4039
rect 950 3967 1140 4005
rect 950 3933 956 3967
rect 990 3933 1028 3967
rect 1062 3966 1140 3967
rect 1062 3933 1100 3966
rect 950 3932 1100 3933
rect 1134 3932 1140 3966
rect 950 3894 1140 3932
rect 950 3860 956 3894
rect 990 3860 1028 3894
rect 1062 3893 1140 3894
rect 1062 3860 1100 3893
rect 950 3859 1100 3860
rect 1134 3859 1140 3893
rect 950 3821 1140 3859
rect 950 3787 956 3821
rect 990 3787 1028 3821
rect 1062 3820 1140 3821
rect 1062 3787 1100 3820
rect 950 3786 1100 3787
rect 1134 3786 1140 3820
rect 950 3748 1140 3786
rect 950 3714 956 3748
rect 990 3714 1028 3748
rect 1062 3747 1140 3748
rect 1062 3714 1100 3747
rect 950 3713 1100 3714
rect 1134 3713 1140 3747
rect 950 3675 1140 3713
rect 950 3641 956 3675
rect 990 3641 1028 3675
rect 1062 3674 1140 3675
rect 1062 3641 1100 3674
rect 950 3640 1100 3641
rect 1134 3640 1140 3674
rect 950 3602 1140 3640
rect 950 3568 956 3602
rect 990 3568 1028 3602
rect 1062 3601 1140 3602
rect 1062 3568 1100 3601
rect 950 3567 1100 3568
rect 1134 3567 1140 3601
rect 950 3529 1140 3567
rect 950 3495 956 3529
rect 990 3495 1028 3529
rect 1062 3528 1140 3529
rect 1062 3495 1100 3528
rect 950 3494 1100 3495
rect 1134 3494 1140 3528
rect 950 3456 1140 3494
rect 950 3422 956 3456
rect 990 3422 1028 3456
rect 1062 3455 1140 3456
rect 1062 3422 1100 3455
rect 950 3421 1100 3422
rect 1134 3421 1140 3455
rect 950 3383 1140 3421
rect 950 3349 956 3383
rect 990 3349 1028 3383
rect 1062 3382 1140 3383
rect 1062 3349 1100 3382
rect 950 3348 1100 3349
rect 1134 3348 1140 3382
rect 950 3310 1140 3348
rect 950 3276 956 3310
rect 990 3276 1028 3310
rect 1062 3309 1140 3310
rect 1062 3276 1100 3309
rect 950 3275 1100 3276
rect 1134 3275 1140 3309
rect 950 3237 1140 3275
rect 950 3203 956 3237
rect 990 3203 1028 3237
rect 1062 3236 1140 3237
rect 1062 3203 1100 3236
rect 950 3202 1100 3203
rect 1134 3202 1140 3236
rect 950 3164 1140 3202
rect 950 3130 956 3164
rect 990 3130 1028 3164
rect 1062 3163 1140 3164
rect 1062 3130 1100 3163
rect 950 3129 1100 3130
rect 1134 3129 1140 3163
rect 950 3091 1140 3129
rect 950 3057 956 3091
rect 990 3057 1028 3091
rect 1062 3090 1140 3091
rect 1062 3057 1100 3090
rect 950 3056 1100 3057
rect 1134 3056 1140 3090
rect 950 3018 1140 3056
rect 950 2984 956 3018
rect 990 2984 1028 3018
rect 1062 3017 1140 3018
rect 1062 2984 1100 3017
rect 950 2983 1100 2984
rect 1134 2983 1140 3017
rect 950 2945 1140 2983
rect 950 2911 956 2945
rect 990 2911 1028 2945
rect 1062 2944 1140 2945
rect 1062 2911 1100 2944
rect 950 2910 1100 2911
rect 1134 2910 1140 2944
rect 950 2872 1140 2910
rect 950 2838 956 2872
rect 990 2838 1028 2872
rect 1062 2871 1140 2872
rect 1062 2838 1100 2871
rect 950 2837 1100 2838
rect 1134 2837 1140 2871
rect 950 2799 1140 2837
rect 950 2765 956 2799
rect 990 2765 1028 2799
rect 1062 2798 1140 2799
rect 1062 2765 1100 2798
rect 950 2764 1100 2765
rect 1134 2764 1140 2798
rect 950 2726 1140 2764
rect 950 2692 956 2726
rect 990 2692 1028 2726
rect 1062 2725 1140 2726
rect 1062 2692 1100 2725
rect 950 2691 1100 2692
rect 1134 2691 1140 2725
rect 950 2653 1140 2691
rect 950 2619 956 2653
rect 990 2619 1028 2653
rect 1062 2652 1140 2653
rect 1062 2619 1100 2652
rect 950 2618 1100 2619
rect 1134 2618 1140 2652
rect 950 2580 1140 2618
rect 950 2546 956 2580
rect 990 2546 1028 2580
rect 1062 2579 1140 2580
rect 1062 2546 1100 2579
rect 950 2545 1100 2546
rect 1134 2545 1140 2579
rect 950 2507 1140 2545
rect 950 2473 956 2507
rect 990 2473 1028 2507
rect 1062 2506 1140 2507
rect 1062 2473 1100 2506
rect 950 2472 1100 2473
rect 1134 2472 1140 2506
rect 950 2434 1140 2472
rect 950 2400 956 2434
rect 990 2400 1028 2434
rect 1062 2433 1140 2434
rect 1062 2400 1100 2433
rect 950 2399 1100 2400
rect 1134 2399 1140 2433
rect 950 2361 1140 2399
rect 950 2327 956 2361
rect 990 2327 1028 2361
rect 1062 2360 1140 2361
rect 1062 2327 1100 2360
rect 950 2326 1100 2327
rect 1134 2326 1140 2360
rect 950 2288 1140 2326
rect 950 2254 956 2288
rect 990 2254 1028 2288
rect 1062 2287 1140 2288
rect 1062 2254 1100 2287
rect 950 2253 1100 2254
rect 1134 2253 1140 2287
rect 950 2215 1140 2253
rect 950 2181 956 2215
rect 990 2181 1028 2215
rect 1062 2214 1140 2215
rect 1062 2181 1100 2214
rect 950 2180 1100 2181
rect 1134 2180 1140 2214
rect 950 2142 1140 2180
rect 950 2108 956 2142
rect 990 2108 1028 2142
rect 1062 2141 1140 2142
rect 1062 2108 1100 2141
rect 950 2107 1100 2108
rect 1134 2107 1140 2141
rect 950 2069 1140 2107
rect 950 2035 956 2069
rect 990 2035 1028 2069
rect 1062 2068 1140 2069
rect 1062 2035 1100 2068
rect 950 2034 1100 2035
rect 1134 2034 1140 2068
rect 950 1996 1140 2034
rect 950 1962 956 1996
rect 990 1962 1028 1996
rect 1062 1995 1140 1996
rect 1062 1962 1100 1995
rect 950 1961 1100 1962
rect 1134 1961 1140 1995
rect 950 1923 1140 1961
rect 950 1889 956 1923
rect 990 1889 1028 1923
rect 1062 1922 1140 1923
rect 1062 1889 1100 1922
rect 950 1888 1100 1889
rect 1134 1888 1140 1922
rect 950 1850 1140 1888
rect 950 1816 956 1850
rect 990 1816 1028 1850
rect 1062 1849 1140 1850
rect 1062 1816 1100 1849
rect 950 1815 1100 1816
rect 1134 1815 1140 1849
rect 950 1777 1140 1815
rect 950 1743 956 1777
rect 990 1743 1028 1777
rect 1062 1776 1140 1777
rect 1062 1743 1100 1776
rect 950 1742 1100 1743
rect 1134 1742 1140 1776
rect 25873 7353 26063 7391
rect 25873 7319 25879 7353
rect 25913 7351 26063 7353
rect 25913 7319 25951 7351
rect 25873 7317 25951 7319
rect 25985 7317 26023 7351
rect 26057 7317 26063 7351
rect 25873 7279 26063 7317
rect 25873 7245 25879 7279
rect 25913 7277 26063 7279
rect 25913 7245 25951 7277
rect 25873 7243 25951 7245
rect 25985 7243 26023 7277
rect 26057 7243 26063 7277
rect 25873 7205 26063 7243
rect 25873 7171 25879 7205
rect 25913 7204 26063 7205
rect 25913 7171 25951 7204
rect 25873 7170 25951 7171
rect 25985 7170 26023 7204
rect 26057 7170 26063 7204
rect 25873 7131 26063 7170
rect 25873 7097 25879 7131
rect 25913 7097 25951 7131
rect 25985 7097 26023 7131
rect 26057 7097 26063 7131
rect 25873 7021 26063 7097
rect 25873 6987 25879 7021
rect 25913 6987 25951 7021
rect 25985 6987 26023 7021
rect 26057 6987 26063 7021
rect 25873 6948 26063 6987
rect 25873 6914 25879 6948
rect 25913 6914 25951 6948
rect 25985 6914 26023 6948
rect 26057 6914 26063 6948
rect 25873 6875 26063 6914
rect 25873 6841 25879 6875
rect 25913 6841 25951 6875
rect 25985 6841 26023 6875
rect 26057 6841 26063 6875
rect 25873 6802 26063 6841
rect 25873 6768 25879 6802
rect 25913 6768 25951 6802
rect 25985 6768 26023 6802
rect 26057 6768 26063 6802
rect 25873 6729 26063 6768
rect 25873 6695 25879 6729
rect 25913 6695 25951 6729
rect 25985 6695 26023 6729
rect 26057 6695 26063 6729
rect 25873 6656 26063 6695
rect 25873 6622 25879 6656
rect 25913 6622 25951 6656
rect 25985 6622 26023 6656
rect 26057 6622 26063 6656
rect 25873 6583 26063 6622
rect 25873 6549 25879 6583
rect 25913 6549 25951 6583
rect 25985 6549 26023 6583
rect 26057 6549 26063 6583
rect 25873 6510 26063 6549
rect 25873 6476 25879 6510
rect 25913 6476 25951 6510
rect 25985 6476 26023 6510
rect 26057 6476 26063 6510
rect 25873 6437 26063 6476
rect 25873 6403 25879 6437
rect 25913 6403 25951 6437
rect 25985 6403 26023 6437
rect 26057 6403 26063 6437
rect 25873 6364 26063 6403
rect 25873 6330 25879 6364
rect 25913 6330 25951 6364
rect 25985 6330 26023 6364
rect 26057 6330 26063 6364
rect 25873 6291 26063 6330
rect 25873 6257 25879 6291
rect 25913 6257 25951 6291
rect 25985 6257 26023 6291
rect 26057 6257 26063 6291
rect 25873 6218 26063 6257
rect 25873 6184 25879 6218
rect 25913 6184 25951 6218
rect 25985 6184 26023 6218
rect 26057 6184 26063 6218
rect 25873 6145 26063 6184
rect 25873 6111 25879 6145
rect 25913 6111 25951 6145
rect 25985 6111 26023 6145
rect 26057 6111 26063 6145
rect 25873 6072 26063 6111
rect 25873 6038 25879 6072
rect 25913 6038 25951 6072
rect 25985 6038 26023 6072
rect 26057 6038 26063 6072
rect 25873 5999 26063 6038
rect 25873 5965 25879 5999
rect 25913 5965 25951 5999
rect 25985 5965 26023 5999
rect 26057 5965 26063 5999
rect 25873 5926 26063 5965
rect 25873 5892 25879 5926
rect 25913 5892 25951 5926
rect 25985 5892 26023 5926
rect 26057 5892 26063 5926
rect 25873 5853 26063 5892
rect 25873 5819 25879 5853
rect 25913 5819 25951 5853
rect 25985 5819 26023 5853
rect 26057 5819 26063 5853
rect 25873 5780 26063 5819
rect 25873 5746 25879 5780
rect 25913 5746 25951 5780
rect 25985 5746 26023 5780
rect 26057 5746 26063 5780
rect 25873 5707 26063 5746
rect 25873 5673 25879 5707
rect 25913 5673 25951 5707
rect 25985 5673 26023 5707
rect 26057 5673 26063 5707
rect 25873 5634 26063 5673
rect 25873 5600 25879 5634
rect 25913 5600 25951 5634
rect 25985 5600 26023 5634
rect 26057 5600 26063 5634
rect 25873 5561 26063 5600
rect 25873 5527 25879 5561
rect 25913 5527 25951 5561
rect 25985 5527 26023 5561
rect 26057 5527 26063 5561
rect 25873 5488 26063 5527
rect 25873 5454 25879 5488
rect 25913 5454 25951 5488
rect 25985 5454 26023 5488
rect 26057 5454 26063 5488
rect 25873 5415 26063 5454
rect 25873 5381 25879 5415
rect 25913 5381 25951 5415
rect 25985 5381 26023 5415
rect 26057 5381 26063 5415
rect 25873 5342 26063 5381
rect 25873 5308 25879 5342
rect 25913 5308 25951 5342
rect 25985 5308 26023 5342
rect 26057 5308 26063 5342
rect 25873 5269 26063 5308
rect 25873 5235 25879 5269
rect 25913 5235 25951 5269
rect 25985 5235 26023 5269
rect 26057 5235 26063 5269
rect 25873 5196 26063 5235
rect 25873 5162 25879 5196
rect 25913 5162 25951 5196
rect 25985 5162 26023 5196
rect 26057 5162 26063 5196
rect 25873 5123 26063 5162
rect 25873 5089 25879 5123
rect 25913 5089 25951 5123
rect 25985 5089 26023 5123
rect 26057 5089 26063 5123
rect 25873 5050 26063 5089
rect 25873 5016 25879 5050
rect 25913 5016 25951 5050
rect 25985 5016 26023 5050
rect 26057 5016 26063 5050
rect 25873 4977 26063 5016
rect 25873 4943 25879 4977
rect 25913 4943 25951 4977
rect 25985 4943 26023 4977
rect 26057 4943 26063 4977
rect 25873 4904 26063 4943
rect 25873 4870 25879 4904
rect 25913 4870 25951 4904
rect 25985 4870 26023 4904
rect 26057 4870 26063 4904
rect 25873 4831 26063 4870
rect 25873 4797 25879 4831
rect 25913 4797 25951 4831
rect 25985 4797 26023 4831
rect 26057 4797 26063 4831
rect 25873 4758 26063 4797
rect 25873 4724 25879 4758
rect 25913 4724 25951 4758
rect 25985 4724 26023 4758
rect 26057 4724 26063 4758
rect 25873 4685 26063 4724
rect 25873 4651 25879 4685
rect 25913 4651 25951 4685
rect 25985 4651 26023 4685
rect 26057 4651 26063 4685
rect 25873 4612 26063 4651
rect 25873 4578 25879 4612
rect 25913 4578 25951 4612
rect 25985 4578 26023 4612
rect 26057 4578 26063 4612
rect 25873 4539 26063 4578
rect 25873 4505 25879 4539
rect 25913 4505 25951 4539
rect 25985 4505 26023 4539
rect 26057 4505 26063 4539
rect 25873 4466 26063 4505
rect 25873 4432 25879 4466
rect 25913 4432 25951 4466
rect 25985 4432 26023 4466
rect 26057 4432 26063 4466
rect 25873 4393 26063 4432
rect 25873 4359 25879 4393
rect 25913 4359 25951 4393
rect 25985 4359 26023 4393
rect 26057 4359 26063 4393
rect 25873 4320 26063 4359
rect 25873 4286 25879 4320
rect 25913 4286 25951 4320
rect 25985 4286 26023 4320
rect 26057 4286 26063 4320
rect 25873 4247 26063 4286
rect 25873 4213 25879 4247
rect 25913 4213 25951 4247
rect 25985 4213 26023 4247
rect 26057 4213 26063 4247
rect 25873 4174 26063 4213
rect 25873 4140 25879 4174
rect 25913 4140 25951 4174
rect 25985 4140 26023 4174
rect 26057 4140 26063 4174
rect 25873 4101 26063 4140
rect 25873 4067 25879 4101
rect 25913 4067 25951 4101
rect 25985 4067 26023 4101
rect 26057 4067 26063 4101
rect 25873 4028 26063 4067
rect 25873 3994 25879 4028
rect 25913 3994 25951 4028
rect 25985 3994 26023 4028
rect 26057 3994 26063 4028
rect 25873 3955 26063 3994
rect 25873 3921 25879 3955
rect 25913 3921 25951 3955
rect 25985 3921 26023 3955
rect 26057 3921 26063 3955
rect 25873 3882 26063 3921
rect 25873 3848 25879 3882
rect 25913 3848 25951 3882
rect 25985 3848 26023 3882
rect 26057 3848 26063 3882
rect 25873 3809 26063 3848
rect 25873 3775 25879 3809
rect 25913 3775 25951 3809
rect 25985 3775 26023 3809
rect 26057 3775 26063 3809
rect 25873 3736 26063 3775
rect 25873 3702 25879 3736
rect 25913 3702 25951 3736
rect 25985 3702 26023 3736
rect 26057 3702 26063 3736
rect 25873 3663 26063 3702
rect 25873 3629 25879 3663
rect 25913 3629 25951 3663
rect 25985 3629 26023 3663
rect 26057 3629 26063 3663
rect 25873 3590 26063 3629
rect 25873 3556 25879 3590
rect 25913 3556 25951 3590
rect 25985 3556 26023 3590
rect 26057 3556 26063 3590
rect 25873 3517 26063 3556
rect 25873 3483 25879 3517
rect 25913 3483 25951 3517
rect 25985 3483 26023 3517
rect 26057 3483 26063 3517
rect 25873 3444 26063 3483
rect 25873 3410 25879 3444
rect 25913 3410 25951 3444
rect 25985 3410 26023 3444
rect 26057 3410 26063 3444
rect 25873 3371 26063 3410
rect 25873 3337 25879 3371
rect 25913 3337 25951 3371
rect 25985 3337 26023 3371
rect 26057 3337 26063 3371
rect 25873 3298 26063 3337
rect 25873 3264 25879 3298
rect 25913 3264 25951 3298
rect 25985 3264 26023 3298
rect 26057 3264 26063 3298
rect 25873 3225 26063 3264
rect 25873 3191 25879 3225
rect 25913 3191 25951 3225
rect 25985 3191 26023 3225
rect 26057 3191 26063 3225
rect 25873 3152 26063 3191
rect 25873 3118 25879 3152
rect 25913 3118 25951 3152
rect 25985 3118 26023 3152
rect 26057 3118 26063 3152
rect 25873 3079 26063 3118
rect 25873 3045 25879 3079
rect 25913 3045 25951 3079
rect 25985 3045 26023 3079
rect 26057 3045 26063 3079
rect 25873 3006 26063 3045
rect 25873 2972 25879 3006
rect 25913 2972 25951 3006
rect 25985 2972 26023 3006
rect 26057 2972 26063 3006
rect 25873 2933 26063 2972
rect 25873 2899 25879 2933
rect 25913 2899 25951 2933
rect 25985 2899 26023 2933
rect 26057 2899 26063 2933
rect 25873 2860 26063 2899
rect 25873 2826 25879 2860
rect 25913 2826 25951 2860
rect 25985 2826 26023 2860
rect 26057 2826 26063 2860
rect 25873 2787 26063 2826
rect 25873 2753 25879 2787
rect 25913 2753 25951 2787
rect 25985 2753 26023 2787
rect 26057 2753 26063 2787
rect 25873 2714 26063 2753
rect 25873 2680 25879 2714
rect 25913 2680 25951 2714
rect 25985 2680 26023 2714
rect 26057 2680 26063 2714
rect 25873 2641 26063 2680
rect 25873 2607 25879 2641
rect 25913 2607 25951 2641
rect 25985 2607 26023 2641
rect 26057 2607 26063 2641
rect 25873 2568 26063 2607
rect 25873 2534 25879 2568
rect 25913 2534 25951 2568
rect 25985 2534 26023 2568
rect 26057 2534 26063 2568
rect 25873 2495 26063 2534
rect 950 1709 1140 1742
tri 1140 1709 1200 1769 sw
tri 25813 1709 25873 1769 se
rect 25873 1709 25879 2495
rect 950 1704 25879 1709
rect 950 1670 956 1704
rect 990 1670 1028 1704
rect 1062 1703 25879 1704
rect 1062 1670 1100 1703
rect 950 1631 1100 1670
rect 25110 1669 25149 1703
rect 25183 1669 25222 1703
rect 25256 1669 25295 1703
rect 25329 1669 25368 1703
rect 25402 1669 25441 1703
rect 25475 1669 25514 1703
rect 25548 1669 25587 1703
rect 25621 1669 25660 1703
rect 25694 1669 25733 1703
rect 25767 1669 25806 1703
rect 25840 1669 25879 1703
rect 25110 1631 25951 1669
rect 950 1597 956 1631
rect 990 1597 1028 1631
rect 950 1525 1028 1597
rect 25182 1597 25221 1631
rect 25255 1597 25294 1631
rect 25328 1597 25367 1631
rect 25401 1597 25440 1631
rect 25474 1597 25513 1631
rect 25547 1597 25586 1631
rect 25620 1597 25659 1631
rect 25693 1597 25732 1631
rect 25766 1597 25805 1631
rect 25839 1597 25878 1631
rect 25912 1597 25951 1631
rect 26057 1597 26063 2495
rect 25182 1559 26063 1597
rect 25182 1525 25221 1559
rect 25255 1525 25294 1559
rect 25328 1525 25367 1559
rect 25401 1525 25440 1559
rect 25474 1525 25513 1559
rect 25547 1525 25586 1559
rect 25620 1525 25659 1559
rect 25693 1525 25732 1559
rect 25766 1525 25805 1559
rect 25839 1525 25878 1559
rect 25912 1525 25951 1559
rect 25985 1525 26063 1559
rect 950 1519 26063 1525
rect 26271 7705 26277 7739
rect 26311 7737 26461 7739
rect 26311 7705 26349 7737
rect 26271 7703 26349 7705
rect 26383 7703 26421 7737
rect 26455 7703 26461 7737
rect 26271 7665 26461 7703
rect 26271 7631 26277 7665
rect 26311 7663 26461 7665
rect 26311 7631 26349 7663
rect 26271 7629 26349 7631
rect 26383 7629 26421 7663
rect 26455 7629 26461 7663
rect 26271 7591 26461 7629
rect 26271 7557 26277 7591
rect 26311 7590 26461 7591
rect 26311 7557 26349 7590
rect 26271 7556 26349 7557
rect 26383 7556 26421 7590
rect 26455 7556 26461 7590
rect 26271 7517 26461 7556
rect 26271 7483 26277 7517
rect 26311 7483 26349 7517
rect 26383 7483 26421 7517
rect 26455 7483 26461 7517
rect 26271 7407 26461 7483
rect 26271 7373 26277 7407
rect 26311 7373 26349 7407
rect 26383 7373 26421 7407
rect 26455 7373 26461 7407
rect 26271 7334 26461 7373
rect 26271 7300 26277 7334
rect 26311 7300 26349 7334
rect 26383 7300 26421 7334
rect 26455 7300 26461 7334
rect 26271 7261 26461 7300
rect 26271 7227 26277 7261
rect 26311 7227 26349 7261
rect 26383 7227 26421 7261
rect 26455 7227 26461 7261
rect 26271 7188 26461 7227
rect 26271 7154 26277 7188
rect 26311 7154 26349 7188
rect 26383 7154 26421 7188
rect 26455 7154 26461 7188
rect 26271 7115 26461 7154
rect 26271 7081 26277 7115
rect 26311 7081 26349 7115
rect 26383 7081 26421 7115
rect 26455 7081 26461 7115
rect 26271 7042 26461 7081
rect 564 1476 570 1510
rect 604 1476 642 1510
rect 676 1509 754 1510
rect 676 1476 714 1509
rect 564 1475 714 1476
rect 748 1475 754 1509
rect 564 1437 754 1475
rect 564 1403 570 1437
rect 604 1403 642 1437
rect 676 1436 754 1437
rect 676 1403 714 1436
rect 564 1402 714 1403
rect 748 1402 754 1436
rect 564 1364 754 1402
rect 564 1330 570 1364
rect 604 1330 642 1364
rect 676 1363 754 1364
rect 676 1330 714 1363
rect 564 1329 714 1330
rect 748 1329 754 1363
rect 564 1291 754 1329
rect 564 1257 570 1291
rect 604 1257 642 1291
rect 676 1290 754 1291
rect 676 1257 714 1290
rect 564 1256 714 1257
rect 748 1256 754 1290
rect 564 1218 754 1256
rect 564 1184 570 1218
rect 604 1184 642 1218
rect 676 1217 754 1218
rect 676 1184 714 1217
rect 564 1183 714 1184
rect 748 1183 754 1217
rect 564 1145 754 1183
rect 564 1111 570 1145
rect 604 1111 642 1145
rect 676 1144 754 1145
rect 676 1111 714 1144
rect 564 1110 714 1111
rect 748 1110 754 1144
rect 564 1072 754 1110
rect 564 1038 570 1072
rect 604 1038 642 1072
rect 676 1071 754 1072
rect 676 1038 714 1071
rect 564 1037 714 1038
rect 748 1037 754 1071
rect 564 999 754 1037
rect 564 965 570 999
rect 604 965 642 999
rect 676 998 754 999
rect 676 965 714 998
rect 564 964 714 965
rect 748 964 754 998
rect 564 926 754 964
rect 564 892 570 926
rect 604 892 642 926
rect 676 925 754 926
rect 676 892 714 925
rect 564 891 714 892
rect 748 891 754 925
rect 564 853 754 891
rect 564 819 570 853
rect 604 819 642 853
rect 676 852 754 853
rect 676 819 714 852
rect 564 818 714 819
rect 748 818 754 852
rect 564 780 754 818
rect 564 746 570 780
rect 604 746 642 780
rect 676 779 754 780
rect 676 746 714 779
rect 564 745 714 746
rect 748 745 754 779
rect 564 712 754 745
tri 754 712 833 791 sw
tri 26211 712 26271 772 se
rect 26271 712 26277 7042
rect 564 707 26277 712
rect 564 673 570 707
rect 604 673 642 707
rect 676 706 26277 707
rect 676 673 714 706
rect 564 634 714 673
rect 26092 672 26131 706
rect 26165 672 26204 706
rect 26238 672 26277 706
rect 26092 634 26349 672
rect 564 600 570 634
rect 604 600 642 634
rect 564 528 642 600
rect 26164 600 26203 634
rect 26237 600 26276 634
rect 26310 600 26349 634
rect 26455 600 26461 7042
rect 26164 562 26461 600
rect 26164 528 26203 562
rect 26237 528 26276 562
rect 26310 528 26349 562
rect 26383 528 26461 562
rect 564 522 26461 528
rect 26674 8099 26680 8133
rect 26714 8099 26752 8133
rect 26786 8099 26824 8133
rect 26858 8099 26864 8133
rect 26674 8054 26864 8099
rect 26674 8020 26680 8054
rect 26714 8020 26752 8054
rect 26786 8020 26824 8054
rect 26858 8020 26864 8054
rect 26674 7975 26864 8020
rect 26674 7941 26680 7975
rect 26714 7941 26752 7975
rect 26786 7941 26824 7975
rect 26858 7941 26864 7975
rect 26674 7896 26864 7941
rect 26674 7862 26680 7896
rect 26714 7862 26752 7896
rect 26786 7862 26824 7896
rect 26858 7862 26864 7896
rect 26674 7786 26864 7862
rect 26674 7752 26680 7786
rect 26714 7752 26752 7786
rect 26786 7752 26824 7786
rect 26858 7752 26864 7786
rect 26674 7713 26864 7752
rect 26674 7679 26680 7713
rect 26714 7679 26752 7713
rect 26786 7679 26824 7713
rect 26858 7679 26864 7713
rect 26674 7640 26864 7679
rect 26674 7606 26680 7640
rect 26714 7606 26752 7640
rect 26786 7606 26824 7640
rect 26858 7606 26864 7640
rect 26674 7567 26864 7606
rect 26674 7533 26680 7567
rect 26714 7533 26752 7567
rect 26786 7533 26824 7567
rect 26858 7533 26864 7567
rect 26674 7494 26864 7533
rect 116 481 306 519
rect 116 447 122 481
rect 156 447 194 481
rect 228 480 306 481
rect 228 447 266 480
rect 116 446 266 447
rect 300 446 306 480
rect 116 408 306 446
rect 116 374 122 408
rect 156 374 194 408
rect 228 407 306 408
rect 228 374 266 407
rect 116 373 266 374
rect 300 373 306 407
rect 116 340 306 373
tri 306 340 366 400 sw
tri 26614 340 26674 400 se
rect 26674 340 26680 7494
rect 116 335 26680 340
rect 116 301 122 335
rect 156 301 194 335
rect 228 334 26680 335
rect 228 301 266 334
rect 116 262 266 301
rect 22548 300 22587 334
rect 22621 300 22660 334
rect 22694 300 22733 334
rect 22767 300 22806 334
rect 22840 300 22879 334
rect 22913 300 22952 334
rect 22986 300 23025 334
rect 23059 300 23098 334
rect 23132 300 23171 334
rect 23205 300 23244 334
rect 23278 300 23317 334
rect 23351 300 23390 334
rect 23424 300 23463 334
rect 23497 300 23536 334
rect 23570 300 23609 334
rect 23643 300 23682 334
rect 23716 300 23755 334
rect 23789 300 23828 334
rect 23862 300 23901 334
rect 23935 300 23974 334
rect 24008 300 24047 334
rect 24081 300 24120 334
rect 24154 300 24193 334
rect 24227 300 24266 334
rect 24300 300 24339 334
rect 24373 300 24412 334
rect 24446 300 24485 334
rect 24519 300 24558 334
rect 24592 300 24631 334
rect 24665 300 24704 334
rect 24738 300 24777 334
rect 24811 300 24850 334
rect 24884 300 24923 334
rect 24957 300 24996 334
rect 25030 300 25069 334
rect 25103 300 25142 334
rect 25176 300 25215 334
rect 25249 300 25288 334
rect 25322 300 25361 334
rect 25395 300 25434 334
rect 25468 300 25507 334
rect 25541 300 25580 334
rect 25614 300 25653 334
rect 25687 300 25726 334
rect 25760 300 25799 334
rect 25833 300 25872 334
rect 25906 300 25945 334
rect 25979 300 26018 334
rect 26052 300 26091 334
rect 26125 300 26164 334
rect 26198 300 26237 334
rect 26271 300 26310 334
rect 26344 300 26383 334
rect 26417 300 26456 334
rect 26490 300 26529 334
rect 26563 300 26602 334
rect 26636 300 26680 334
rect 22548 262 26680 300
rect 116 228 122 262
rect 156 228 194 262
rect 116 156 194 228
rect 22548 228 22587 262
rect 22621 228 22660 262
rect 22694 228 22733 262
rect 22767 228 22806 262
rect 22840 228 22879 262
rect 22913 228 22952 262
rect 22986 228 23025 262
rect 23059 228 23098 262
rect 23132 228 23171 262
rect 23205 228 23244 262
rect 23278 228 23317 262
rect 23351 228 23390 262
rect 23424 228 23463 262
rect 23497 228 23536 262
rect 23570 228 23609 262
rect 23643 228 23682 262
rect 23716 228 23755 262
rect 23789 228 23828 262
rect 23862 228 23901 262
rect 23935 228 23974 262
rect 24008 228 24047 262
rect 24081 228 24120 262
rect 24154 228 24193 262
rect 24227 228 24266 262
rect 24300 228 24339 262
rect 24373 228 24412 262
rect 24446 228 24485 262
rect 24519 228 24558 262
rect 24592 228 24631 262
rect 24665 228 24704 262
rect 24738 228 24777 262
rect 24811 228 24850 262
rect 24884 228 24923 262
rect 24957 228 24996 262
rect 25030 228 25069 262
rect 25103 228 25142 262
rect 25176 228 25215 262
rect 25249 228 25288 262
rect 25322 228 25361 262
rect 25395 228 25434 262
rect 25468 228 25507 262
rect 25541 228 25580 262
rect 25614 228 25653 262
rect 25687 228 25726 262
rect 25760 228 25799 262
rect 25833 228 25872 262
rect 25906 228 25945 262
rect 25979 228 26018 262
rect 26052 228 26091 262
rect 26125 228 26164 262
rect 26198 228 26237 262
rect 26271 228 26310 262
rect 26344 228 26383 262
rect 26417 228 26456 262
rect 26490 228 26529 262
rect 26563 228 26602 262
rect 26636 228 26680 262
rect 22548 190 26680 228
rect 22548 156 22587 190
rect 22621 156 22660 190
rect 22694 156 22733 190
rect 22767 156 22806 190
rect 22840 156 22879 190
rect 22913 156 22952 190
rect 22986 156 23025 190
rect 23059 156 23098 190
rect 23132 156 23171 190
rect 23205 156 23244 190
rect 23278 156 23317 190
rect 23351 156 23390 190
rect 23424 156 23463 190
rect 23497 156 23536 190
rect 23570 156 23609 190
rect 23643 156 23682 190
rect 23716 156 23755 190
rect 23789 156 23828 190
rect 23862 156 23901 190
rect 23935 156 23974 190
rect 24008 156 24047 190
rect 24081 156 24120 190
rect 24154 156 24193 190
rect 24227 156 24266 190
rect 24300 156 24339 190
rect 24373 156 24412 190
rect 24446 156 24485 190
rect 24519 156 24558 190
rect 24592 156 24631 190
rect 24665 156 24704 190
rect 24738 156 24777 190
rect 24811 156 24850 190
rect 24884 156 24923 190
rect 24957 156 24996 190
rect 25030 156 25069 190
rect 25103 156 25142 190
rect 25176 156 25215 190
rect 25249 156 25288 190
rect 25322 156 25361 190
rect 25395 156 25434 190
rect 25468 156 25507 190
rect 25541 156 25580 190
rect 25614 156 25653 190
rect 25687 156 25726 190
rect 25760 156 25799 190
rect 25833 156 25872 190
rect 25906 156 25945 190
rect 25979 156 26018 190
rect 26052 156 26091 190
rect 26125 156 26164 190
rect 26198 156 26237 190
rect 26271 156 26310 190
rect 26344 156 26383 190
rect 26417 156 26456 190
rect 26490 156 26529 190
rect 26563 156 26602 190
rect 26636 188 26680 190
rect 26858 188 26864 7494
rect 26636 156 26864 188
rect 116 150 26864 156
<< properties >>
string GDS_END 35259966
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 34175442
<< end >>
