/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield.model.spice