magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 0 2 5 6 6 DRAIN
port 1 nsew
rlabel rotate s 4 8 4 8 6 GATE
port 2 nsew
rlabel rotate s 4 0 4 0 8 GATE
port 2 nsew
rlabel rotate s 3 8 4 8 6 GATE
port 2 nsew
rlabel rotate s 3 0 4 0 8 GATE
port 2 nsew
rlabel rotate s 3 8 3 8 6 GATE
port 2 nsew
rlabel rotate s 3 0 3 0 8 GATE
port 2 nsew
rlabel rotate s 3 8 3 8 6 GATE
port 2 nsew
rlabel rotate s 3 0 3 0 8 GATE
port 2 nsew
rlabel rotate s 2 8 2 8 6 GATE
port 2 nsew
rlabel rotate s 2 0 2 0 8 GATE
port 2 nsew
rlabel rotate s 2 8 2 8 6 GATE
port 2 nsew
rlabel rotate s 2 0 2 0 8 GATE
port 2 nsew
rlabel rotate s 2 8 2 8 6 GATE
port 2 nsew
rlabel rotate s 2 0 2 0 8 GATE
port 2 nsew
rlabel rotate s 1 8 1 8 6 GATE
port 2 nsew
rlabel rotate s 1 0 1 0 8 GATE
port 2 nsew
rlabel  s 1 8 4 8 6 GATE
port 2 nsew
rlabel  s 1 0 4 0 8 GATE
port 2 nsew
rlabel  s 1 8 4 8 6 GATE
port 2 nsew
rlabel  s 1 0 4 0 8 GATE
port 2 nsew
rlabel  s 0 6 5 7 6 SOURCE
port 3 nsew
rlabel  s 0 1 5 2 6 SOURCE
port 3 nsew
rlabel  s 0 1 0 7 4 SUBSTRATE
port 4 nsew
rlabel  s 5 1 5 7 6 SUBSTRATE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 5 8
string LEFview TRUE
<< end >>
