/home/nataraj/projects/designmyic/cad/pdk/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice