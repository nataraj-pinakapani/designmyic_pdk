magic
tech minimum
magscale 1 2
timestamp 1644097982
<< labels >>
rlabel  s 4 9 4 12 6 GATE
port 1 nsew
rlabel rotate s 4 9 4 9 6 GATE
port 1 nsew
rlabel rotate s 4 9 4 9 6 GATE
port 1 nsew
rlabel � s 3 9 5 9 6 GATE
port 1 nsew
rlabel  s 5 0 7 0 8 NWELLRING
port 2 nsew
rlabel  s 0 0 1 0 2 NWELLRING
port 2 nsew
rlabel  s 5 0 7 1 8 NWELLRING
port 2 nsew
rlabel  s 7 1 7 1 6 NWELLRING
port 2 nsew
rlabel  s 7 1 8 11 6 NWELLRING
port 2 nsew
rlabel  s 7 11 8 11 6 NWELLRING
port 2 nsew
rlabel  s 7 11 8 11 6 NWELLRING
port 2 nsew
rlabel  s 0 0 1 11 4 NWELLRING
port 2 nsew
rlabel  s 6 11 7 11 6 NWELLRING
port 2 nsew
rlabel  s 1 11 1 11 6 NWELLRING
port 2 nsew
rlabel  s 4 11 7 12 6 NWELLRING
port 2 nsew
rlabel  s 1 11 3 12 6 NWELLRING
port 2 nsew
rlabel rotate s 6 1 6 1 6 NWELLRING
port 2 nsew
rlabel rotate s 6 1 6 1 6 NWELLRING
port 2 nsew
rlabel rotate s 6 1 6 1 6 NWELLRING
port 2 nsew
rlabel rotate s 7 1 7 2 6 NWELLRING
port 2 nsew
rlabel rotate s 7 2 7 2 6 NWELLRING
port 2 nsew
rlabel rotate s 7 2 7 2 6 NWELLRING
port 2 nsew
rlabel rotate s 7 2 7 3 6 NWELLRING
port 2 nsew
rlabel rotate s 7 3 7 3 6 NWELLRING
port 2 nsew
rlabel rotate s 7 3 7 3 6 NWELLRING
port 2 nsew
rlabel rotate s 7 4 7 4 6 NWELLRING
port 2 nsew
rlabel rotate s 7 4 7 4 6 NWELLRING
port 2 nsew
rlabel rotate s 7 4 7 4 6 NWELLRING
port 2 nsew
rlabel rotate s 7 5 7 5 6 NWELLRING
port 2 nsew
rlabel rotate s 7 5 7 5 6 NWELLRING
port 2 nsew
rlabel rotate s 7 5 7 5 6 NWELLRING
port 2 nsew
rlabel rotate s 7 6 7 6 6 NWELLRING
port 2 nsew
rlabel rotate s 7 6 7 6 6 NWELLRING
port 2 nsew
rlabel rotate s 7 6 7 7 6 NWELLRING
port 2 nsew
rlabel rotate s 7 7 7 7 6 NWELLRING
port 2 nsew
rlabel rotate s 7 7 7 7 6 NWELLRING
port 2 nsew
rlabel rotate s 7 7 7 8 6 NWELLRING
port 2 nsew
rlabel rotate s 7 8 7 8 6 NWELLRING
port 2 nsew
rlabel rotate s 7 8 7 8 6 NWELLRING
port 2 nsew
rlabel rotate s 7 9 7 9 6 NWELLRING
port 2 nsew
rlabel rotate s 7 9 7 9 6 NWELLRING
port 2 nsew
rlabel rotate s 7 9 7 9 6 NWELLRING
port 2 nsew
rlabel rotate s 7 10 7 10 6 NWELLRING
port 2 nsew
rlabel rotate s 7 10 7 10 6 NWELLRING
port 2 nsew
rlabel rotate s 1 1 1 2 6 NWELLRING
port 2 nsew
rlabel rotate s 1 2 1 2 6 NWELLRING
port 2 nsew
rlabel rotate s 1 2 1 2 6 NWELLRING
port 2 nsew
rlabel rotate s 1 2 1 3 6 NWELLRING
port 2 nsew
rlabel rotate s 1 3 1 3 6 NWELLRING
port 2 nsew
rlabel rotate s 1 3 1 3 6 NWELLRING
port 2 nsew
rlabel rotate s 1 4 1 4 6 NWELLRING
port 2 nsew
rlabel rotate s 1 4 1 4 6 NWELLRING
port 2 nsew
rlabel rotate s 1 4 1 4 6 NWELLRING
port 2 nsew
rlabel rotate s 1 5 1 5 6 NWELLRING
port 2 nsew
rlabel rotate s 1 5 1 5 6 NWELLRING
port 2 nsew
rlabel rotate s 1 5 1 5 6 NWELLRING
port 2 nsew
rlabel rotate s 1 6 1 6 6 NWELLRING
port 2 nsew
rlabel rotate s 1 6 1 6 6 NWELLRING
port 2 nsew
rlabel rotate s 1 6 1 7 6 NWELLRING
port 2 nsew
rlabel rotate s 1 7 1 7 6 NWELLRING
port 2 nsew
rlabel rotate s 1 7 1 7 6 NWELLRING
port 2 nsew
rlabel rotate s 1 7 1 8 6 NWELLRING
port 2 nsew
rlabel rotate s 1 8 1 8 6 NWELLRING
port 2 nsew
rlabel rotate s 1 8 1 8 6 NWELLRING
port 2 nsew
rlabel rotate s 1 9 1 9 6 NWELLRING
port 2 nsew
rlabel rotate s 1 9 1 9 6 NWELLRING
port 2 nsew
rlabel rotate s 1 9 1 9 6 NWELLRING
port 2 nsew
rlabel rotate s 1 10 1 10 6 NWELLRING
port 2 nsew
rlabel rotate s 1 10 1 10 6 NWELLRING
port 2 nsew
rlabel rotate s 6 11 6 12 6 NWELLRING
port 2 nsew
rlabel rotate s 6 11 6 12 6 NWELLRING
port 2 nsew
rlabel rotate s 6 11 6 12 6 NWELLRING
port 2 nsew
rlabel rotate s 5 11 5 12 6 NWELLRING
port 2 nsew
rlabel rotate s 5 11 5 12 6 NWELLRING
port 2 nsew
rlabel rotate s 3 11 3 12 6 NWELLRING
port 2 nsew
rlabel rotate s 3 11 3 12 6 NWELLRING
port 2 nsew
rlabel rotate s 2 11 2 12 6 NWELLRING
port 2 nsew
rlabel rotate s 2 11 2 12 6 NWELLRING
port 2 nsew
rlabel rotate s 2 11 2 12 6 NWELLRING
port 2 nsew
rlabel � s 0 0 8 1 8 NWELLRING
port 2 nsew
rlabel � s 7 1 8 11 6 NWELLRING
port 2 nsew
rlabel � s 0 1 1 11 4 NWELLRING
port 2 nsew
rlabel � s 0 11 8 12 6 NWELLRING
port 2 nsew
rlabel dark_red s 0 0 8 1 8 NWELLRING
port 2 nsew
rlabel dark_red s 7 1 8 11 6 NWELLRING
port 2 nsew
rlabel dark_red s 0 1 1 11 4 NWELLRING
port 2 nsew
rlabel dark_red s 0 11 8 12 6 NWELLRING
port 2 nsew
rlabel  s 3 0 4 9 6 VGND
port 3 nsew ground default
rlabel rotate s 3 4 3 4 6 VGND
port 3 nsew ground default
rlabel rotate s 3 4 3 4 6 VGND
port 3 nsew ground default
rlabel rotate s 3 5 3 5 6 VGND
port 3 nsew ground default
rlabel rotate s 3 5 3 5 6 VGND
port 3 nsew ground default
rlabel rotate s 3 5 3 5 6 VGND
port 3 nsew ground default
rlabel rotate s 3 6 3 6 6 VGND
port 3 nsew ground default
rlabel rotate s 3 6 3 6 6 VGND
port 3 nsew ground default
rlabel rotate s 3 6 3 6 6 VGND
port 3 nsew ground default
rlabel rotate s 3 7 3 7 6 VGND
port 3 nsew ground default
rlabel rotate s 3 7 3 7 6 VGND
port 3 nsew ground default
rlabel rotate s 3 7 3 8 6 VGND
port 3 nsew ground default
rlabel rotate s 3 8 3 8 6 VGND
port 3 nsew ground default
rlabel � s 3 3 4 9 6 VGND
port 3 nsew ground default
rlabel  s 2 0 3 0 8 NBODY
port 4 nsew
rlabel  s 5 2 6 9 6 NBODY
port 4 nsew
rlabel  s 5 9 6 10 6 NBODY
port 4 nsew
rlabel  s 2 0 3 10 6 NBODY
port 4 nsew
rlabel  s 4 10 6 10 6 NBODY
port 4 nsew
rlabel  s 4 10 6 10 6 NBODY
port 4 nsew
rlabel  s 2 10 3 10 6 NBODY
port 4 nsew
rlabel  s 2 10 3 10 6 NBODY
port 4 nsew
rlabel rotate s 6 2 6 2 6 NBODY
port 4 nsew
rlabel rotate s 2 2 2 2 6 NBODY
port 4 nsew
rlabel rotate s 6 2 6 3 6 NBODY
port 4 nsew
rlabel rotate s 6 3 6 3 6 NBODY
port 4 nsew
rlabel rotate s 6 3 6 3 6 NBODY
port 4 nsew
rlabel rotate s 6 3 6 4 6 NBODY
port 4 nsew
rlabel rotate s 6 4 6 4 6 NBODY
port 4 nsew
rlabel rotate s 6 4 6 4 6 NBODY
port 4 nsew
rlabel rotate s 6 5 6 5 6 NBODY
port 4 nsew
rlabel rotate s 6 5 6 5 6 NBODY
port 4 nsew
rlabel rotate s 6 5 6 5 6 NBODY
port 4 nsew
rlabel rotate s 6 6 6 6 6 NBODY
port 4 nsew
rlabel rotate s 6 6 6 6 6 NBODY
port 4 nsew
rlabel rotate s 6 6 6 6 6 NBODY
port 4 nsew
rlabel rotate s 6 7 6 7 6 NBODY
port 4 nsew
rlabel rotate s 6 7 6 7 6 NBODY
port 4 nsew
rlabel rotate s 6 7 6 8 6 NBODY
port 4 nsew
rlabel rotate s 6 8 6 8 6 NBODY
port 4 nsew
rlabel rotate s 6 8 6 8 6 NBODY
port 4 nsew
rlabel rotate s 6 8 6 9 6 NBODY
port 4 nsew
rlabel rotate s 6 9 6 9 6 NBODY
port 4 nsew
rlabel rotate s 2 2 2 3 6 NBODY
port 4 nsew
rlabel rotate s 2 3 2 3 6 NBODY
port 4 nsew
rlabel rotate s 2 3 2 3 6 NBODY
port 4 nsew
rlabel rotate s 2 3 2 4 6 NBODY
port 4 nsew
rlabel rotate s 2 4 2 4 6 NBODY
port 4 nsew
rlabel rotate s 2 4 2 4 6 NBODY
port 4 nsew
rlabel rotate s 2 5 2 5 6 NBODY
port 4 nsew
rlabel rotate s 2 5 2 5 6 NBODY
port 4 nsew
rlabel rotate s 2 5 2 5 6 NBODY
port 4 nsew
rlabel rotate s 2 6 2 6 6 NBODY
port 4 nsew
rlabel rotate s 2 6 2 6 6 NBODY
port 4 nsew
rlabel rotate s 2 6 2 6 6 NBODY
port 4 nsew
rlabel rotate s 2 7 2 7 6 NBODY
port 4 nsew
rlabel rotate s 2 7 2 7 6 NBODY
port 4 nsew
rlabel rotate s 2 7 2 8 6 NBODY
port 4 nsew
rlabel rotate s 2 8 2 8 6 NBODY
port 4 nsew
rlabel rotate s 2 8 2 8 6 NBODY
port 4 nsew
rlabel rotate s 2 8 2 9 6 NBODY
port 4 nsew
rlabel rotate s 2 9 2 9 6 NBODY
port 4 nsew
rlabel rotate s 5 10 6 10 6 NBODY
port 4 nsew
rlabel rotate s 5 10 5 10 6 NBODY
port 4 nsew
rlabel rotate s 5 10 5 10 6 NBODY
port 4 nsew
rlabel rotate s 3 10 3 10 6 NBODY
port 4 nsew
rlabel rotate s 3 10 3 10 6 NBODY
port 4 nsew
rlabel rotate s 2 10 2 10 6 NBODY
port 4 nsew
rlabel � s 2 2 6 2 6 NBODY
port 4 nsew
rlabel � s 5 2 6 10 6 NBODY
port 4 nsew
rlabel � s 2 2 2 10 6 NBODY
port 4 nsew
rlabel � s 2 10 6 10 6 NBODY
port 4 nsew
rlabel metal_blue s 2 2 6 10 6 NBODY
port 4 nsew
rlabel  s 4 0 5 9 6 IN
port 5 nsew
rlabel rotate s 5 4 5 4 6 IN
port 5 nsew
rlabel rotate s 5 4 5 4 6 IN
port 5 nsew
rlabel rotate s 5 5 5 5 6 IN
port 5 nsew
rlabel rotate s 5 5 5 5 6 IN
port 5 nsew
rlabel rotate s 5 5 5 5 6 IN
port 5 nsew
rlabel rotate s 5 6 5 6 6 IN
port 5 nsew
rlabel rotate s 5 6 5 6 6 IN
port 5 nsew
rlabel rotate s 5 6 5 6 6 IN
port 5 nsew
rlabel rotate s 5 7 5 7 6 IN
port 5 nsew
rlabel rotate s 5 7 5 7 6 IN
port 5 nsew
rlabel rotate s 5 7 5 8 6 IN
port 5 nsew
rlabel rotate s 5 8 5 8 6 IN
port 5 nsew
rlabel � s 4 3 5 9 6 IN
port 5 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 8 12
string LEFview TRUE
<< end >>
