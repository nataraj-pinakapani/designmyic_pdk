magic
tech sky130B
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 24 21 1256 203
rect 25 -17 59 21
<< scnmos >>
rect 102 47 132 177
rect 186 47 216 177
rect 276 47 306 177
rect 360 47 390 177
rect 552 47 582 177
rect 636 47 666 177
rect 728 47 758 177
rect 812 47 842 177
rect 896 47 926 177
rect 980 47 1010 177
rect 1064 47 1094 177
rect 1148 47 1178 177
<< scpmoshvt >>
rect 102 297 132 497
rect 186 297 216 497
rect 276 297 306 497
rect 360 297 390 497
rect 444 297 474 497
rect 532 297 562 497
rect 728 297 758 497
rect 812 297 842 497
rect 896 297 926 497
rect 980 297 1010 497
rect 1064 297 1094 497
rect 1148 297 1178 497
<< ndiff >>
rect 50 93 102 177
rect 50 59 58 93
rect 92 59 102 93
rect 50 47 102 59
rect 132 161 186 177
rect 132 127 142 161
rect 176 127 186 161
rect 132 47 186 127
rect 216 89 276 177
rect 216 55 229 89
rect 263 55 276 89
rect 216 47 276 55
rect 306 161 360 177
rect 306 127 316 161
rect 350 127 360 161
rect 306 47 360 127
rect 390 161 442 177
rect 390 127 400 161
rect 434 127 442 161
rect 390 93 442 127
rect 390 59 400 93
rect 434 59 442 93
rect 390 47 442 59
rect 496 89 552 177
rect 496 55 508 89
rect 542 55 552 89
rect 496 47 552 55
rect 582 169 636 177
rect 582 135 592 169
rect 626 135 636 169
rect 582 47 636 135
rect 666 129 728 177
rect 666 95 678 129
rect 712 95 728 129
rect 666 47 728 95
rect 758 89 812 177
rect 758 55 768 89
rect 802 55 812 89
rect 758 47 812 55
rect 842 129 896 177
rect 842 95 852 129
rect 886 95 896 129
rect 842 47 896 95
rect 926 89 980 177
rect 926 55 936 89
rect 970 55 980 89
rect 926 47 980 55
rect 1010 129 1064 177
rect 1010 95 1020 129
rect 1054 95 1064 129
rect 1010 47 1064 95
rect 1094 89 1148 177
rect 1094 55 1104 89
rect 1138 55 1148 89
rect 1094 47 1148 55
rect 1178 129 1230 177
rect 1178 95 1188 129
rect 1222 95 1230 129
rect 1178 47 1230 95
<< pdiff >>
rect 50 485 102 497
rect 50 451 58 485
rect 92 451 102 485
rect 50 417 102 451
rect 50 383 58 417
rect 92 383 102 417
rect 50 297 102 383
rect 132 448 186 497
rect 132 414 142 448
rect 176 414 186 448
rect 132 380 186 414
rect 132 346 142 380
rect 176 346 186 380
rect 132 297 186 346
rect 216 489 276 497
rect 216 455 229 489
rect 263 455 276 489
rect 216 421 276 455
rect 216 387 229 421
rect 263 387 276 421
rect 216 297 276 387
rect 306 448 360 497
rect 306 414 316 448
rect 350 414 360 448
rect 306 380 360 414
rect 306 346 316 380
rect 350 346 360 380
rect 306 297 360 346
rect 390 489 444 497
rect 390 455 400 489
rect 434 455 444 489
rect 390 421 444 455
rect 390 387 400 421
rect 434 387 444 421
rect 390 353 444 387
rect 390 319 400 353
rect 434 319 444 353
rect 390 297 444 319
rect 474 448 532 497
rect 474 414 488 448
rect 522 414 532 448
rect 474 380 532 414
rect 474 346 488 380
rect 522 346 532 380
rect 474 297 532 346
rect 562 489 618 497
rect 562 455 572 489
rect 606 455 618 489
rect 562 297 618 455
rect 672 340 728 497
rect 672 306 684 340
rect 718 306 728 340
rect 672 297 728 306
rect 758 489 812 497
rect 758 455 768 489
rect 802 455 812 489
rect 758 421 812 455
rect 758 387 768 421
rect 802 387 812 421
rect 758 297 812 387
rect 842 448 896 497
rect 842 414 852 448
rect 886 414 896 448
rect 842 380 896 414
rect 842 346 852 380
rect 886 346 896 380
rect 842 297 896 346
rect 926 424 980 497
rect 926 390 936 424
rect 970 390 980 424
rect 926 297 980 390
rect 1010 489 1064 497
rect 1010 455 1020 489
rect 1054 455 1064 489
rect 1010 297 1064 455
rect 1094 424 1148 497
rect 1094 390 1104 424
rect 1138 390 1148 424
rect 1094 297 1148 390
rect 1178 448 1230 497
rect 1178 414 1188 448
rect 1222 414 1230 448
rect 1178 297 1230 414
<< ndiffc >>
rect 58 59 92 93
rect 142 127 176 161
rect 229 55 263 89
rect 316 127 350 161
rect 400 127 434 161
rect 400 59 434 93
rect 508 55 542 89
rect 592 135 626 169
rect 678 95 712 129
rect 768 55 802 89
rect 852 95 886 129
rect 936 55 970 89
rect 1020 95 1054 129
rect 1104 55 1138 89
rect 1188 95 1222 129
<< pdiffc >>
rect 58 451 92 485
rect 58 383 92 417
rect 142 414 176 448
rect 142 346 176 380
rect 229 455 263 489
rect 229 387 263 421
rect 316 414 350 448
rect 316 346 350 380
rect 400 455 434 489
rect 400 387 434 421
rect 400 319 434 353
rect 488 414 522 448
rect 488 346 522 380
rect 572 455 606 489
rect 684 306 718 340
rect 768 455 802 489
rect 768 387 802 421
rect 852 414 886 448
rect 852 346 886 380
rect 936 390 970 424
rect 1020 455 1054 489
rect 1104 390 1138 424
rect 1188 414 1222 448
<< poly >>
rect 102 497 132 523
rect 186 497 216 523
rect 276 497 306 523
rect 360 497 390 523
rect 444 497 474 523
rect 532 497 562 523
rect 728 497 758 523
rect 812 497 842 523
rect 896 497 926 523
rect 980 497 1010 523
rect 1064 497 1094 523
rect 1148 497 1178 523
rect 102 259 132 297
rect 186 259 216 297
rect 276 259 306 297
rect 360 259 390 297
rect 102 249 390 259
rect 102 215 204 249
rect 238 215 272 249
rect 306 215 340 249
rect 374 215 390 249
rect 102 205 390 215
rect 444 259 474 297
rect 532 259 562 297
rect 728 259 758 297
rect 812 259 842 297
rect 896 265 926 297
rect 444 249 666 259
rect 444 215 608 249
rect 642 215 666 249
rect 444 205 666 215
rect 102 177 132 205
rect 186 177 216 205
rect 276 177 306 205
rect 360 177 390 205
rect 552 177 582 205
rect 636 177 666 205
rect 728 249 842 259
rect 728 215 769 249
rect 803 215 842 249
rect 728 205 842 215
rect 728 177 758 205
rect 812 177 842 205
rect 884 249 938 265
rect 884 215 894 249
rect 928 215 938 249
rect 884 199 938 215
rect 980 259 1010 297
rect 1064 259 1094 297
rect 980 249 1094 259
rect 980 215 1044 249
rect 1078 215 1094 249
rect 980 205 1094 215
rect 896 177 926 199
rect 980 177 1010 205
rect 1064 177 1094 205
rect 1148 259 1178 297
rect 1148 249 1214 259
rect 1148 215 1164 249
rect 1198 215 1214 249
rect 1148 205 1214 215
rect 1148 177 1178 205
rect 102 21 132 47
rect 186 21 216 47
rect 276 21 306 47
rect 360 21 390 47
rect 552 21 582 47
rect 636 21 666 47
rect 728 21 758 47
rect 812 21 842 47
rect 896 21 926 47
rect 980 21 1010 47
rect 1064 21 1094 47
rect 1148 21 1178 47
<< polycont >>
rect 204 215 238 249
rect 272 215 306 249
rect 340 215 374 249
rect 608 215 642 249
rect 769 215 803 249
rect 894 215 928 249
rect 1044 215 1078 249
rect 1164 215 1198 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 485 102 527
rect 17 451 58 485
rect 92 451 102 485
rect 17 417 102 451
rect 17 383 58 417
rect 92 383 102 417
rect 17 367 102 383
rect 136 448 179 493
rect 136 414 142 448
rect 176 414 179 448
rect 136 380 179 414
rect 136 346 142 380
rect 176 346 179 380
rect 213 489 279 527
rect 213 455 229 489
rect 263 455 279 489
rect 213 421 279 455
rect 213 387 229 421
rect 263 387 279 421
rect 213 367 279 387
rect 313 448 350 493
rect 313 414 316 448
rect 313 380 350 414
rect 136 333 179 346
rect 313 346 316 380
rect 313 333 350 346
rect 17 292 350 333
rect 384 489 450 527
rect 384 455 400 489
rect 434 455 450 489
rect 384 421 450 455
rect 384 387 400 421
rect 434 387 450 421
rect 384 353 450 387
rect 384 319 400 353
rect 434 319 450 353
rect 384 292 450 319
rect 488 448 522 493
rect 556 489 622 527
rect 556 455 572 489
rect 606 455 622 489
rect 556 448 622 455
rect 752 489 818 493
rect 752 455 768 489
rect 802 455 818 489
rect 752 421 818 455
rect 752 414 768 421
rect 488 387 768 414
rect 802 387 818 421
rect 488 380 818 387
rect 522 374 818 380
rect 852 459 902 493
rect 852 448 857 459
rect 891 425 902 459
rect 886 414 902 425
rect 852 380 902 414
rect 17 177 147 292
rect 488 258 522 346
rect 886 346 902 380
rect 936 424 970 493
rect 1004 489 1070 527
rect 1004 455 1020 489
rect 1054 455 1070 489
rect 1004 448 1070 455
rect 1104 424 1144 493
rect 970 390 1104 414
rect 1138 390 1144 424
rect 936 374 1144 390
rect 1178 459 1271 493
rect 1178 448 1225 459
rect 1178 414 1188 448
rect 1222 425 1225 448
rect 1259 425 1271 459
rect 1222 414 1271 425
rect 1178 374 1271 414
rect 852 340 902 346
rect 181 249 522 258
rect 181 215 204 249
rect 238 215 272 249
rect 306 215 340 249
rect 374 215 522 249
rect 181 211 522 215
rect 556 271 630 339
rect 664 306 684 340
rect 718 306 902 340
rect 936 306 1271 340
rect 936 272 994 306
rect 556 249 715 271
rect 556 215 608 249
rect 642 215 715 249
rect 556 211 715 215
rect 753 249 819 272
rect 753 215 769 249
rect 803 215 819 249
rect 753 211 819 215
rect 853 249 994 272
rect 853 215 894 249
rect 928 215 994 249
rect 853 211 994 215
rect 1028 249 1094 272
rect 1028 215 1044 249
rect 1078 215 1094 249
rect 1028 211 1094 215
rect 1128 249 1271 306
rect 1128 215 1164 249
rect 1198 215 1271 249
rect 1128 211 1271 215
rect 488 177 522 211
rect 17 161 353 177
rect 17 143 142 161
rect 136 127 142 143
rect 176 131 316 161
rect 176 127 179 131
rect 17 93 102 109
rect 17 59 58 93
rect 92 59 102 93
rect 17 17 102 59
rect 136 51 179 127
rect 313 127 316 131
rect 350 127 353 161
rect 213 89 279 97
rect 213 55 229 89
rect 263 55 279 89
rect 213 17 279 55
rect 313 51 353 127
rect 387 161 450 177
rect 387 127 400 161
rect 434 127 450 161
rect 488 169 642 177
rect 488 135 592 169
rect 626 135 642 169
rect 488 127 642 135
rect 676 129 1271 177
rect 387 93 450 127
rect 676 95 678 129
rect 712 127 852 129
rect 712 95 714 127
rect 676 93 714 95
rect 387 59 400 93
rect 434 59 450 93
rect 387 17 450 59
rect 488 89 714 93
rect 886 127 1020 129
rect 488 55 508 89
rect 542 55 714 89
rect 488 51 714 55
rect 752 55 768 89
rect 802 55 818 89
rect 752 17 818 55
rect 852 51 886 95
rect 1054 127 1188 129
rect 920 55 936 89
rect 970 55 986 89
rect 920 17 986 55
rect 1020 51 1054 95
rect 1222 95 1271 129
rect 1088 55 1104 89
rect 1138 55 1154 89
rect 1088 17 1154 55
rect 1188 51 1271 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 857 448 891 459
rect 857 425 886 448
rect 886 425 891 448
rect 1225 425 1259 459
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 845 459 903 465
rect 845 425 857 459
rect 891 456 903 459
rect 1213 459 1271 465
rect 1213 456 1225 459
rect 891 428 1225 456
rect 891 425 903 428
rect 845 419 903 425
rect 1213 425 1225 428
rect 1259 425 1271 459
rect 1213 419 1271 425
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 25 153 59 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 113 153 147 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 113 221 147 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 25 221 59 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 25 289 59 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 113 289 147 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 577 289 611 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 577 221 611 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 669 221 703 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 949 289 983 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1133 289 1167 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1225 289 1259 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel metal1 s 25 -17 59 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 25 527 59 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 25 527 59 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 25 -17 59 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o31a_4
rlabel metal1 s 0 -48 1288 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 1423826
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_sc_hd/sky130_fd_sc_hd.gds
string GDS_START 1412714
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 6.440 2.720 
<< end >>
