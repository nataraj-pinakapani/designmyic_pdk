* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******* SkyWater sky130 model library *********
.subckt sky130_all_dummy
.ends
* Typical corner (tt)
.lib tt
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl tt

* Slow-Fast corner (sf)
.lib sf
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/sf.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/sf/specialized_cells.spice"
.endl sf

* Fast-Fast corner (ff)
.lib ff
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/ff.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/ff/specialized_cells.spice"
.endl ff

* Slow-Slow corner (ss)
.lib ss
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/ss.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/ss/specialized_cells.spice"
.endl ss

* Fast-Slow corner (fs)
.lib fs
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/fs.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/fs/specialized_cells.spice"
.endl fs

* Low-Low corner (ll)
.lib ll
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_low__cap_low.spice"
.include "r+c/res_low__cap_low__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl ll

* High-High corner (hh)
.lib hh
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_high__cap_high.spice"
.include "r+c/res_high__cap_high__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl hh

* High-Low corner (hl)
.lib hl
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_high__cap_low.spice"
.include "r+c/res_high__cap_low__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl hl

* Low-High corner (lh)
.lib lh
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_low__cap_high.spice"
.include "r+c/res_low__cap_high__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl lh

* Typical corner with mismatch (tt_mm)
.lib tt_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl tt_mm

* Slow-Fast corner with mismatch (sf_mm)
.lib sf_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/sf.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/sf/specialized_cells.spice"
.endl sf_mm

* Fast-Fast corner with mismatch (ff_mm)
.lib ff_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/ff.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/ff/specialized_cells.spice"
.endl ff_mm

* Slow-Slow corner with mismatch (ss_mm)
.lib ss_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/ss.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/ss/specialized_cells.spice"
.endl ss_mm

* Fast-Slow corner with mismatch (fs_mm)
.lib fs_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/fs.spice"
* Resistor/Capacitor
.include "r+c/res_typical__cap_typical.spice"
.include "r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "corners/fs/specialized_cells.spice"
.endl fs_mm

* Low-Low corner with mismatch (ll_mm)
.lib ll_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_low__cap_low.spice"
.include "r+c/res_low__cap_low__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl ll_mm

* High-High corner with mismatch (hh_mm)
.lib hh_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_high__cap_high.spice"
.include "r+c/res_high__cap_high__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl hh_mm

* High-Low corner with mismatch (hl_mm)
.lib hl_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_high__cap_low.spice"
.include "r+c/res_high__cap_low__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl hl_mm

* Low-High corner with mismatch (lh_mm)
.lib lh_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "corners/tt.spice"
* Resistor/Capacitor
.include "r+c/res_low__cap_high.spice"
.include "r+c/res_low__cap_high__lin.spice"
* Special cells
.include "corners/tt/specialized_cells.spice"
.endl lh_mm

* Monte Carlo process variation

.lib mc

.param mc_mm_switch=0
.param mc_pr_switch=1

.include "parameters/critical.spice"
.include "parameters/montecarlo.spice"

.endl mc
