magic
tech minimum
magscale 1 2
timestamp 1644097874
<< labels >>
rlabel  s 17 8 17 15 6 C0
port 1 nsew
rlabel  s 17 0 17 8 6 C0
port 1 nsew
rlabel  s 15 12 16 15 6 C0
port 1 nsew
rlabel  s 15 8 16 11 6 C0
port 1 nsew
rlabel  s 15 4 16 8 6 C0
port 1 nsew
rlabel  s 15 0 16 3 6 C0
port 1 nsew
rlabel  s 14 12 14 15 6 C0
port 1 nsew
rlabel  s 14 8 14 11 6 C0
port 1 nsew
rlabel  s 14 4 14 8 6 C0
port 1 nsew
rlabel  s 14 0 14 3 6 C0
port 1 nsew
rlabel  s 12 12 13 15 6 C0
port 1 nsew
rlabel  s 12 8 13 11 6 C0
port 1 nsew
rlabel  s 12 4 13 8 6 C0
port 1 nsew
rlabel  s 12 0 13 3 6 C0
port 1 nsew
rlabel  s 11 12 11 15 6 C0
port 1 nsew
rlabel  s 11 8 11 11 6 C0
port 1 nsew
rlabel  s 11 4 11 8 6 C0
port 1 nsew
rlabel  s 11 0 11 3 6 C0
port 1 nsew
rlabel  s 10 12 10 15 6 C0
port 1 nsew
rlabel  s 10 8 10 11 6 C0
port 1 nsew
rlabel  s 10 4 10 8 6 C0
port 1 nsew
rlabel  s 10 0 10 3 6 C0
port 1 nsew
rlabel  s 8 8 9 15 6 C0
port 1 nsew
rlabel  s 8 0 9 8 6 C0
port 1 nsew
rlabel  s 7 12 7 15 6 C0
port 1 nsew
rlabel  s 7 8 7 11 6 C0
port 1 nsew
rlabel  s 7 4 7 8 6 C0
port 1 nsew
rlabel  s 7 0 7 3 6 C0
port 1 nsew
rlabel  s 5 12 6 15 6 C0
port 1 nsew
rlabel  s 5 8 6 11 6 C0
port 1 nsew
rlabel  s 5 4 6 8 6 C0
port 1 nsew
rlabel  s 5 0 6 3 6 C0
port 1 nsew
rlabel  s 4 12 4 15 6 C0
port 1 nsew
rlabel  s 4 8 4 11 6 C0
port 1 nsew
rlabel  s 4 4 4 8 6 C0
port 1 nsew
rlabel  s 4 0 4 3 6 C0
port 1 nsew
rlabel  s 3 12 3 15 6 C0
port 1 nsew
rlabel  s 3 8 3 11 6 C0
port 1 nsew
rlabel  s 3 4 3 8 6 C0
port 1 nsew
rlabel  s 3 0 3 3 6 C0
port 1 nsew
rlabel  s 1 12 2 15 6 C0
port 1 nsew
rlabel  s 1 8 2 11 6 C0
port 1 nsew
rlabel  s 1 4 2 8 6 C0
port 1 nsew
rlabel  s 1 0 2 3 6 C0
port 1 nsew
rlabel  s 0 15 17 15 6 C0
port 1 nsew
rlabel  s 0 8 0 15 4 C0
port 1 nsew
rlabel  s 0 8 17 8 6 C0
port 1 nsew
rlabel  s 0 0 0 8 4 C0
port 1 nsew
rlabel  s 0 0 17 0 8 C0
port 1 nsew
rlabel  s 16 12 16 15 6 C1
port 2 nsew
rlabel  s 16 8 16 11 6 C1
port 2 nsew
rlabel  s 16 4 16 7 6 C1
port 2 nsew
rlabel  s 16 1 16 4 6 C1
port 2 nsew
rlabel  s 14 12 15 15 6 C1
port 2 nsew
rlabel  s 14 8 15 11 6 C1
port 2 nsew
rlabel  s 14 4 15 7 6 C1
port 2 nsew
rlabel  s 14 1 15 4 6 C1
port 2 nsew
rlabel  s 13 12 13 15 6 C1
port 2 nsew
rlabel  s 13 8 13 11 6 C1
port 2 nsew
rlabel  s 13 4 13 7 6 C1
port 2 nsew
rlabel  s 13 1 13 4 6 C1
port 2 nsew
rlabel  s 12 12 12 15 6 C1
port 2 nsew
rlabel  s 12 8 12 11 6 C1
port 2 nsew
rlabel  s 12 4 12 7 6 C1
port 2 nsew
rlabel  s 12 1 12 4 6 C1
port 2 nsew
rlabel  s 10 12 11 15 6 C1
port 2 nsew
rlabel  s 10 8 11 11 6 C1
port 2 nsew
rlabel  s 10 4 11 7 6 C1
port 2 nsew
rlabel  s 10 1 11 4 6 C1
port 2 nsew
rlabel  s 9 12 9 15 6 C1
port 2 nsew
rlabel  s 9 11 16 12 6 C1
port 2 nsew
rlabel  s 9 8 9 11 6 C1
port 2 nsew
rlabel  s 9 4 9 7 6 C1
port 2 nsew
rlabel  s 9 4 16 4 6 C1
port 2 nsew
rlabel  s 9 1 9 4 6 C1
port 2 nsew
rlabel  s 8 12 8 15 6 C1
port 2 nsew
rlabel  s 8 8 8 11 6 C1
port 2 nsew
rlabel  s 8 4 8 7 6 C1
port 2 nsew
rlabel  s 8 1 8 4 6 C1
port 2 nsew
rlabel  s 6 12 7 15 6 C1
port 2 nsew
rlabel  s 6 8 7 11 6 C1
port 2 nsew
rlabel  s 6 4 7 7 6 C1
port 2 nsew
rlabel  s 6 1 7 4 6 C1
port 2 nsew
rlabel  s 5 12 5 15 6 C1
port 2 nsew
rlabel  s 5 8 5 11 6 C1
port 2 nsew
rlabel  s 5 4 5 7 6 C1
port 2 nsew
rlabel  s 5 1 5 4 6 C1
port 2 nsew
rlabel  s 3 12 4 15 6 C1
port 2 nsew
rlabel  s 3 8 4 11 6 C1
port 2 nsew
rlabel  s 3 4 4 7 6 C1
port 2 nsew
rlabel  s 3 1 4 4 6 C1
port 2 nsew
rlabel  s 2 12 2 15 6 C1
port 2 nsew
rlabel  s 2 8 2 11 6 C1
port 2 nsew
rlabel  s 2 4 2 7 6 C1
port 2 nsew
rlabel  s 2 1 2 4 6 C1
port 2 nsew
rlabel  s 1 12 1 15 6 C1
port 2 nsew
rlabel  s 1 11 8 12 6 C1
port 2 nsew
rlabel  s 1 8 1 11 6 C1
port 2 nsew
rlabel  s 1 4 1 7 6 C1
port 2 nsew
rlabel  s 1 4 8 4 6 C1
port 2 nsew
rlabel  s 1 1 1 4 6 C1
port 2 nsew
rlabel r s 0 0 17 15 6 M5
port 3 nsew
rlabel metal_blue s 6 6 6 6 6 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 17 15
string LEFview TRUE
<< end >>
