magic
tech sky130A
magscale 1 2
timestamp 1663361622
<< nwell >>
rect -179 1414 -91 2367
rect -19 2173 195 2273
rect 6101 2173 6352 2273
<< pwell >>
rect 2477 1941 3819 2231
rect 2511 1599 3785 1941
rect 6052 888 6401 891
rect 6043 197 6401 888
rect 6043 159 12124 197
rect 5539 73 12124 159
rect 1314 -282 3711 -94
rect -253 -1098 3711 -282
<< psubdiff >>
rect 2503 2171 2596 2205
rect 2630 2171 2669 2205
rect 2703 2171 2741 2205
rect 2775 2171 2813 2205
rect 2847 2171 2885 2205
rect 2919 2171 2957 2205
rect 2991 2171 3029 2205
rect 3063 2171 3101 2205
rect 3135 2171 3173 2205
rect 3207 2171 3245 2205
rect 3279 2171 3317 2205
rect 3351 2171 3389 2205
rect 3423 2171 3461 2205
rect 3495 2171 3533 2205
rect 3567 2171 3605 2205
rect 3639 2171 3677 2205
rect 3711 2171 3793 2205
rect 2503 2137 3793 2171
rect 2503 2103 2596 2137
rect 2630 2103 2669 2137
rect 2703 2103 2741 2137
rect 2775 2103 2813 2137
rect 2847 2103 2885 2137
rect 2919 2103 2957 2137
rect 2991 2103 3029 2137
rect 3063 2103 3101 2137
rect 3135 2103 3173 2137
rect 3207 2103 3245 2137
rect 3279 2103 3317 2137
rect 3351 2103 3389 2137
rect 3423 2103 3461 2137
rect 3495 2103 3533 2137
rect 3567 2103 3605 2137
rect 3639 2103 3677 2137
rect 3711 2103 3793 2137
rect 2503 2069 3793 2103
rect 2503 2035 2596 2069
rect 2630 2035 2669 2069
rect 2703 2035 2741 2069
rect 2775 2035 2813 2069
rect 2847 2035 2885 2069
rect 2919 2035 2957 2069
rect 2991 2035 3029 2069
rect 3063 2035 3101 2069
rect 3135 2035 3173 2069
rect 3207 2035 3245 2069
rect 3279 2035 3317 2069
rect 3351 2035 3389 2069
rect 3423 2035 3461 2069
rect 3495 2035 3533 2069
rect 3567 2035 3605 2069
rect 3639 2035 3677 2069
rect 3711 2035 3793 2069
rect 2503 2001 3793 2035
rect 2503 1967 2596 2001
rect 2630 1967 2669 2001
rect 2703 1967 2741 2001
rect 2775 1967 2813 2001
rect 2847 1967 2885 2001
rect 2919 1967 2957 2001
rect 2991 1967 3029 2001
rect 3063 1967 3101 2001
rect 3135 1967 3173 2001
rect 3207 1967 3245 2001
rect 3279 1967 3317 2001
rect 3351 1967 3389 2001
rect 3423 1967 3461 2001
rect 3495 1967 3533 2001
rect 3567 1967 3605 2001
rect 3639 1967 3677 2001
rect 3711 1967 3793 2001
rect 2537 1933 3759 1967
rect 2537 1899 2579 1933
rect 2613 1899 2648 1933
rect 2682 1899 2717 1933
rect 2751 1899 2786 1933
rect 2820 1899 2855 1933
rect 2889 1899 2924 1933
rect 2958 1899 2993 1933
rect 3027 1899 3062 1933
rect 3096 1899 3131 1933
rect 3165 1899 3200 1933
rect 3234 1899 3269 1933
rect 3303 1899 3338 1933
rect 3372 1899 3407 1933
rect 3441 1899 3476 1933
rect 3510 1899 3545 1933
rect 3579 1899 3613 1933
rect 3647 1899 3681 1933
rect 3715 1899 3759 1933
rect 2537 1853 3759 1899
rect 2537 1819 2579 1853
rect 2613 1819 2648 1853
rect 2682 1819 2717 1853
rect 2751 1819 2786 1853
rect 2820 1819 2855 1853
rect 2889 1819 2924 1853
rect 2958 1819 2993 1853
rect 3027 1819 3062 1853
rect 3096 1819 3131 1853
rect 3165 1819 3200 1853
rect 3234 1819 3269 1853
rect 3303 1819 3338 1853
rect 3372 1819 3407 1853
rect 3441 1819 3476 1853
rect 3510 1819 3545 1853
rect 3579 1819 3613 1853
rect 3647 1819 3681 1853
rect 3715 1819 3759 1853
rect 2537 1773 3759 1819
rect 2537 1739 2579 1773
rect 2613 1739 2648 1773
rect 2682 1739 2717 1773
rect 2751 1739 2786 1773
rect 2820 1739 2855 1773
rect 2889 1739 2924 1773
rect 2958 1739 2993 1773
rect 3027 1739 3062 1773
rect 3096 1739 3131 1773
rect 3165 1739 3200 1773
rect 3234 1739 3269 1773
rect 3303 1739 3338 1773
rect 3372 1739 3407 1773
rect 3441 1739 3476 1773
rect 3510 1739 3545 1773
rect 3579 1739 3613 1773
rect 3647 1739 3681 1773
rect 3715 1739 3759 1773
rect 2537 1693 3759 1739
rect 2537 1659 2579 1693
rect 2613 1659 2648 1693
rect 2682 1659 2717 1693
rect 2751 1659 2786 1693
rect 2820 1659 2855 1693
rect 2889 1659 2924 1693
rect 2958 1659 2993 1693
rect 3027 1659 3062 1693
rect 3096 1659 3131 1693
rect 3165 1659 3200 1693
rect 3234 1659 3269 1693
rect 3303 1659 3338 1693
rect 3372 1659 3407 1693
rect 3441 1659 3476 1693
rect 3510 1659 3545 1693
rect 3579 1659 3613 1693
rect 3647 1659 3681 1693
rect 3715 1659 3759 1693
rect 2537 1625 3759 1659
rect 6078 862 6375 865
rect 6069 841 6375 862
rect 6069 195 6102 841
rect 6204 195 6239 841
rect 6341 195 6375 841
rect 6069 171 6375 195
rect 6069 133 12098 171
rect 5565 99 5649 133
rect 5683 99 5934 133
rect 5968 99 6003 133
rect 6037 99 6072 133
rect 6106 99 6141 133
rect 6175 99 6210 133
rect 6244 99 6279 133
rect 6313 99 6348 133
rect 6382 99 6417 133
rect 6451 99 6486 133
rect 6520 99 6555 133
rect 6589 99 6624 133
rect 6658 99 6693 133
rect 6727 99 6762 133
rect 6796 99 6831 133
rect 6865 99 6900 133
rect 6934 99 6969 133
rect 7003 99 7038 133
rect 7072 99 7107 133
rect 7141 99 7176 133
rect 7210 99 7245 133
rect 7279 99 7314 133
rect 7348 99 7383 133
rect 7417 99 7452 133
rect 7486 99 7521 133
rect 7555 99 7590 133
rect 7624 99 7659 133
rect 7693 99 7728 133
rect 7762 99 7797 133
rect 7831 99 7866 133
rect 7900 99 7935 133
rect 7969 99 8004 133
rect 8038 99 8073 133
rect 8107 99 8142 133
rect 8176 99 8211 133
rect 8245 99 8280 133
rect 8314 99 8349 133
rect 8383 99 8418 133
rect 8452 99 8487 133
rect 8521 99 8556 133
rect 8590 99 8625 133
rect 8659 99 8694 133
rect 8728 99 8763 133
rect 8797 99 8832 133
rect 8866 99 8901 133
rect 8935 99 8970 133
rect 9004 99 9039 133
rect 9073 99 9108 133
rect 9142 99 9177 133
rect 9211 99 9246 133
rect 9280 99 9315 133
rect 9349 99 9384 133
rect 9418 99 9453 133
rect 9487 99 9522 133
rect 9556 99 9591 133
rect 9625 99 9660 133
rect 9694 99 9728 133
rect 9762 99 9796 133
rect 9830 99 9864 133
rect 9898 99 9932 133
rect 9966 99 10000 133
rect 10034 99 10068 133
rect 10102 99 10136 133
rect 10170 99 10204 133
rect 10238 99 10272 133
rect 10306 99 10340 133
rect 10374 99 10408 133
rect 10442 99 10476 133
rect 10510 99 10544 133
rect 10578 99 10612 133
rect 10646 99 10680 133
rect 10714 99 10748 133
rect 10782 99 10816 133
rect 10850 99 10884 133
rect 10918 99 10952 133
rect 10986 99 11020 133
rect 11054 99 11088 133
rect 11122 99 11156 133
rect 11190 99 11224 133
rect 11258 99 11292 133
rect 11326 99 11360 133
rect 11394 99 11428 133
rect 11462 99 11496 133
rect 11530 99 11564 133
rect 11598 99 11632 133
rect 11666 99 11700 133
rect 11734 99 11768 133
rect 11802 99 11836 133
rect 11870 99 11904 133
rect 11938 99 11972 133
rect 12006 99 12040 133
rect 12074 99 12098 133
rect 1340 -124 3685 -120
rect 1340 -158 1374 -124
rect 1408 -158 1445 -124
rect 1479 -158 1516 -124
rect 1550 -158 1587 -124
rect 1621 -158 1657 -124
rect 1691 -158 1727 -124
rect 1761 -158 1797 -124
rect 1831 -158 1867 -124
rect 1901 -158 1937 -124
rect 1971 -158 2007 -124
rect 2041 -158 2077 -124
rect 2111 -158 2147 -124
rect 2181 -158 2217 -124
rect 2251 -158 2287 -124
rect 2321 -158 2357 -124
rect 2391 -158 2427 -124
rect 2461 -158 2497 -124
rect 2531 -158 2567 -124
rect 2601 -158 2637 -124
rect 2671 -158 2707 -124
rect 2741 -158 2777 -124
rect 2811 -158 2847 -124
rect 2881 -158 2917 -124
rect 2951 -158 2987 -124
rect 3021 -158 3057 -124
rect 3091 -158 3127 -124
rect 3161 -158 3197 -124
rect 3231 -158 3267 -124
rect 3301 -158 3337 -124
rect 3371 -158 3407 -124
rect 3441 -158 3477 -124
rect 3511 -158 3547 -124
rect 3581 -158 3617 -124
rect 3651 -158 3685 -124
rect 1340 -194 3685 -158
rect 1340 -228 1374 -194
rect 1408 -228 1445 -194
rect 1479 -228 1516 -194
rect 1550 -228 1587 -194
rect 1621 -228 1657 -194
rect 1691 -228 1727 -194
rect 1761 -228 1797 -194
rect 1831 -228 1867 -194
rect 1901 -228 1937 -194
rect 1971 -228 2007 -194
rect 2041 -228 2077 -194
rect 2111 -228 2147 -194
rect 2181 -228 2217 -194
rect 2251 -228 2287 -194
rect 2321 -228 2357 -194
rect 2391 -228 2427 -194
rect 2461 -228 2497 -194
rect 2531 -228 2567 -194
rect 2601 -228 2637 -194
rect 2671 -228 2707 -194
rect 2741 -228 2777 -194
rect 2811 -228 2847 -194
rect 2881 -228 2917 -194
rect 2951 -228 2987 -194
rect 3021 -228 3057 -194
rect 3091 -228 3127 -194
rect 3161 -228 3197 -194
rect 3231 -228 3267 -194
rect 3301 -228 3337 -194
rect 3371 -228 3407 -194
rect 3441 -228 3477 -194
rect 3511 -228 3547 -194
rect 3581 -228 3617 -194
rect 3651 -228 3685 -194
rect 1340 -264 3685 -228
rect 1340 -298 1374 -264
rect 1408 -298 1445 -264
rect 1479 -298 1516 -264
rect 1550 -298 1587 -264
rect 1621 -298 1657 -264
rect 1691 -298 1727 -264
rect 1761 -298 1797 -264
rect 1831 -298 1867 -264
rect 1901 -298 1937 -264
rect 1971 -298 2007 -264
rect 2041 -298 2077 -264
rect 2111 -298 2147 -264
rect 2181 -298 2217 -264
rect 2251 -298 2287 -264
rect 2321 -298 2357 -264
rect 2391 -298 2427 -264
rect 2461 -298 2497 -264
rect 2531 -298 2567 -264
rect 2601 -298 2637 -264
rect 2671 -298 2707 -264
rect 2741 -298 2777 -264
rect 2811 -298 2847 -264
rect 2881 -298 2917 -264
rect 2951 -298 2987 -264
rect 3021 -298 3057 -264
rect 3091 -298 3127 -264
rect 3161 -298 3197 -264
rect 3231 -298 3267 -264
rect 3301 -298 3337 -264
rect 3371 -298 3407 -264
rect 3441 -298 3477 -264
rect 3511 -298 3547 -264
rect 3581 -298 3617 -264
rect 3651 -298 3685 -264
rect 1340 -308 3685 -298
rect -227 -313 3685 -308
rect -227 -347 -193 -313
rect -159 -347 -123 -313
rect -89 -347 -53 -313
rect -19 -347 17 -313
rect 51 -347 87 -313
rect 121 -347 157 -313
rect 191 -347 227 -313
rect 261 -347 297 -313
rect 331 -347 367 -313
rect 401 -347 437 -313
rect 471 -347 507 -313
rect 541 -347 577 -313
rect 611 -347 647 -313
rect 681 -347 717 -313
rect 751 -347 787 -313
rect 821 -347 857 -313
rect 891 -347 927 -313
rect 961 -347 996 -313
rect 1030 -347 1065 -313
rect 1099 -347 1134 -313
rect 1168 -347 1203 -313
rect 1237 -347 1272 -313
rect 1306 -334 3685 -313
rect 1306 -347 1374 -334
rect -227 -368 1374 -347
rect 1408 -368 1445 -334
rect 1479 -368 1516 -334
rect 1550 -368 1587 -334
rect 1621 -368 1657 -334
rect 1691 -368 1727 -334
rect 1761 -368 1797 -334
rect 1831 -368 1867 -334
rect 1901 -368 1937 -334
rect 1971 -368 2007 -334
rect 2041 -368 2077 -334
rect 2111 -368 2147 -334
rect 2181 -368 2217 -334
rect 2251 -368 2287 -334
rect 2321 -368 2357 -334
rect 2391 -368 2427 -334
rect 2461 -368 2497 -334
rect 2531 -368 2567 -334
rect 2601 -368 2637 -334
rect 2671 -368 2707 -334
rect 2741 -368 2777 -334
rect 2811 -368 2847 -334
rect 2881 -368 2917 -334
rect 2951 -368 2987 -334
rect 3021 -368 3057 -334
rect 3091 -368 3127 -334
rect 3161 -368 3197 -334
rect 3231 -368 3267 -334
rect 3301 -368 3337 -334
rect 3371 -368 3407 -334
rect 3441 -368 3477 -334
rect 3511 -368 3547 -334
rect 3581 -368 3617 -334
rect 3651 -368 3685 -334
rect -227 -385 3685 -368
rect -227 -419 -193 -385
rect -159 -419 -123 -385
rect -89 -419 -53 -385
rect -19 -419 17 -385
rect 51 -419 87 -385
rect 121 -419 157 -385
rect 191 -419 227 -385
rect 261 -419 297 -385
rect 331 -419 367 -385
rect 401 -419 437 -385
rect 471 -419 507 -385
rect 541 -419 577 -385
rect 611 -419 647 -385
rect 681 -419 717 -385
rect 751 -419 787 -385
rect 821 -419 857 -385
rect 891 -419 927 -385
rect 961 -419 996 -385
rect 1030 -419 1065 -385
rect 1099 -419 1134 -385
rect 1168 -419 1203 -385
rect 1237 -419 1272 -385
rect 1306 -404 3685 -385
rect 1306 -419 1374 -404
rect -227 -438 1374 -419
rect 1408 -438 1445 -404
rect 1479 -438 1516 -404
rect 1550 -438 1587 -404
rect 1621 -438 1657 -404
rect 1691 -438 1727 -404
rect 1761 -438 1797 -404
rect 1831 -438 1867 -404
rect 1901 -438 1937 -404
rect 1971 -438 2007 -404
rect 2041 -438 2077 -404
rect 2111 -438 2147 -404
rect 2181 -438 2217 -404
rect 2251 -438 2287 -404
rect 2321 -438 2357 -404
rect 2391 -438 2427 -404
rect 2461 -438 2497 -404
rect 2531 -438 2567 -404
rect 2601 -438 2637 -404
rect 2671 -438 2707 -404
rect 2741 -438 2777 -404
rect 2811 -438 2847 -404
rect 2881 -438 2917 -404
rect 2951 -438 2987 -404
rect 3021 -438 3057 -404
rect 3091 -438 3127 -404
rect 3161 -438 3197 -404
rect 3231 -438 3267 -404
rect 3301 -438 3337 -404
rect 3371 -438 3407 -404
rect 3441 -438 3477 -404
rect 3511 -438 3547 -404
rect 3581 -438 3617 -404
rect 3651 -438 3685 -404
rect -227 -457 3685 -438
rect -227 -491 -193 -457
rect -159 -491 -123 -457
rect -89 -491 -53 -457
rect -19 -491 17 -457
rect 51 -491 87 -457
rect 121 -491 157 -457
rect 191 -491 227 -457
rect 261 -491 297 -457
rect 331 -491 367 -457
rect 401 -491 437 -457
rect 471 -491 507 -457
rect 541 -491 577 -457
rect 611 -491 647 -457
rect 681 -491 717 -457
rect 751 -491 787 -457
rect 821 -491 857 -457
rect 891 -491 927 -457
rect 961 -491 996 -457
rect 1030 -491 1065 -457
rect 1099 -491 1134 -457
rect 1168 -491 1203 -457
rect 1237 -491 1272 -457
rect 1306 -474 3685 -457
rect 1306 -491 1374 -474
rect -227 -508 1374 -491
rect 1408 -508 1445 -474
rect 1479 -508 1516 -474
rect 1550 -508 1587 -474
rect 1621 -508 1657 -474
rect 1691 -508 1727 -474
rect 1761 -508 1797 -474
rect 1831 -508 1867 -474
rect 1901 -508 1937 -474
rect 1971 -508 2007 -474
rect 2041 -508 2077 -474
rect 2111 -508 2147 -474
rect 2181 -508 2217 -474
rect 2251 -508 2287 -474
rect 2321 -508 2357 -474
rect 2391 -508 2427 -474
rect 2461 -508 2497 -474
rect 2531 -508 2567 -474
rect 2601 -508 2637 -474
rect 2671 -508 2707 -474
rect 2741 -508 2777 -474
rect 2811 -508 2847 -474
rect 2881 -508 2917 -474
rect 2951 -508 2987 -474
rect 3021 -508 3057 -474
rect 3091 -508 3127 -474
rect 3161 -508 3197 -474
rect 3231 -508 3267 -474
rect 3301 -508 3337 -474
rect 3371 -508 3407 -474
rect 3441 -508 3477 -474
rect 3511 -508 3547 -474
rect 3581 -508 3617 -474
rect 3651 -508 3685 -474
rect -227 -529 3685 -508
rect -227 -563 -193 -529
rect -159 -563 -123 -529
rect -89 -563 -53 -529
rect -19 -563 17 -529
rect 51 -563 87 -529
rect 121 -563 157 -529
rect 191 -563 227 -529
rect 261 -563 297 -529
rect 331 -563 367 -529
rect 401 -563 437 -529
rect 471 -563 507 -529
rect 541 -563 577 -529
rect 611 -563 647 -529
rect 681 -563 717 -529
rect 751 -563 787 -529
rect 821 -563 857 -529
rect 891 -563 927 -529
rect 961 -563 996 -529
rect 1030 -563 1065 -529
rect 1099 -563 1134 -529
rect 1168 -563 1203 -529
rect 1237 -563 1272 -529
rect 1306 -544 3685 -529
rect 1306 -563 1374 -544
rect -227 -578 1374 -563
rect 1408 -578 1445 -544
rect 1479 -578 1516 -544
rect 1550 -578 1587 -544
rect 1621 -578 1657 -544
rect 1691 -578 1727 -544
rect 1761 -578 1797 -544
rect 1831 -578 1867 -544
rect 1901 -578 1937 -544
rect 1971 -578 2007 -544
rect 2041 -578 2077 -544
rect 2111 -578 2147 -544
rect 2181 -578 2217 -544
rect 2251 -578 2287 -544
rect 2321 -578 2357 -544
rect 2391 -578 2427 -544
rect 2461 -578 2497 -544
rect 2531 -578 2567 -544
rect 2601 -578 2637 -544
rect 2671 -578 2707 -544
rect 2741 -578 2777 -544
rect 2811 -578 2847 -544
rect 2881 -578 2917 -544
rect 2951 -578 2987 -544
rect 3021 -578 3057 -544
rect 3091 -578 3127 -544
rect 3161 -578 3197 -544
rect 3231 -578 3267 -544
rect 3301 -578 3337 -544
rect 3371 -578 3407 -544
rect 3441 -578 3477 -544
rect 3511 -578 3547 -544
rect 3581 -578 3617 -544
rect 3651 -578 3685 -544
rect -227 -601 3685 -578
rect -227 -635 -193 -601
rect -159 -635 -123 -601
rect -89 -635 -53 -601
rect -19 -635 17 -601
rect 51 -635 87 -601
rect 121 -635 157 -601
rect 191 -635 227 -601
rect 261 -635 297 -601
rect 331 -635 367 -601
rect 401 -635 437 -601
rect 471 -635 507 -601
rect 541 -635 577 -601
rect 611 -635 647 -601
rect 681 -635 717 -601
rect 751 -635 787 -601
rect 821 -635 857 -601
rect 891 -635 927 -601
rect 961 -635 996 -601
rect 1030 -635 1065 -601
rect 1099 -635 1134 -601
rect 1168 -635 1203 -601
rect 1237 -635 1272 -601
rect 1306 -614 3685 -601
rect 1306 -635 1374 -614
rect -227 -648 1374 -635
rect 1408 -648 1445 -614
rect 1479 -648 1516 -614
rect 1550 -648 1587 -614
rect 1621 -648 1657 -614
rect 1691 -648 1727 -614
rect 1761 -648 1797 -614
rect 1831 -648 1867 -614
rect 1901 -648 1937 -614
rect 1971 -648 2007 -614
rect 2041 -648 2077 -614
rect 2111 -648 2147 -614
rect 2181 -648 2217 -614
rect 2251 -648 2287 -614
rect 2321 -648 2357 -614
rect 2391 -648 2427 -614
rect 2461 -648 2497 -614
rect 2531 -648 2567 -614
rect 2601 -648 2637 -614
rect 2671 -648 2707 -614
rect 2741 -648 2777 -614
rect 2811 -648 2847 -614
rect 2881 -648 2917 -614
rect 2951 -648 2987 -614
rect 3021 -648 3057 -614
rect 3091 -648 3127 -614
rect 3161 -648 3197 -614
rect 3231 -648 3267 -614
rect 3301 -648 3337 -614
rect 3371 -648 3407 -614
rect 3441 -648 3477 -614
rect 3511 -648 3547 -614
rect 3581 -648 3617 -614
rect 3651 -648 3685 -614
rect -227 -673 3685 -648
rect -227 -707 -193 -673
rect -159 -707 -123 -673
rect -89 -707 -53 -673
rect -19 -707 17 -673
rect 51 -707 87 -673
rect 121 -707 157 -673
rect 191 -707 227 -673
rect 261 -707 297 -673
rect 331 -707 367 -673
rect 401 -707 437 -673
rect 471 -707 507 -673
rect 541 -707 577 -673
rect 611 -707 647 -673
rect 681 -707 717 -673
rect 751 -707 787 -673
rect 821 -707 857 -673
rect 891 -707 927 -673
rect 961 -707 996 -673
rect 1030 -707 1065 -673
rect 1099 -707 1134 -673
rect 1168 -707 1203 -673
rect 1237 -707 1272 -673
rect 1306 -684 3685 -673
rect 1306 -707 1374 -684
rect -227 -718 1374 -707
rect 1408 -718 1445 -684
rect 1479 -718 1516 -684
rect 1550 -718 1587 -684
rect 1621 -718 1657 -684
rect 1691 -718 1727 -684
rect 1761 -718 1797 -684
rect 1831 -718 1867 -684
rect 1901 -718 1937 -684
rect 1971 -718 2007 -684
rect 2041 -718 2077 -684
rect 2111 -718 2147 -684
rect 2181 -718 2217 -684
rect 2251 -718 2287 -684
rect 2321 -718 2357 -684
rect 2391 -718 2427 -684
rect 2461 -718 2497 -684
rect 2531 -718 2567 -684
rect 2601 -718 2637 -684
rect 2671 -718 2707 -684
rect 2741 -718 2777 -684
rect 2811 -718 2847 -684
rect 2881 -718 2917 -684
rect 2951 -718 2987 -684
rect 3021 -718 3057 -684
rect 3091 -718 3127 -684
rect 3161 -718 3197 -684
rect 3231 -718 3267 -684
rect 3301 -718 3337 -684
rect 3371 -718 3407 -684
rect 3441 -718 3477 -684
rect 3511 -718 3547 -684
rect 3581 -718 3617 -684
rect 3651 -718 3685 -684
rect -227 -745 3685 -718
rect -227 -779 -193 -745
rect -159 -779 -123 -745
rect -89 -779 -53 -745
rect -19 -779 17 -745
rect 51 -779 87 -745
rect 121 -779 157 -745
rect 191 -779 227 -745
rect 261 -779 297 -745
rect 331 -779 367 -745
rect 401 -779 437 -745
rect 471 -779 507 -745
rect 541 -779 577 -745
rect 611 -779 647 -745
rect 681 -779 717 -745
rect 751 -779 787 -745
rect 821 -779 857 -745
rect 891 -779 927 -745
rect 961 -779 996 -745
rect 1030 -779 1065 -745
rect 1099 -779 1134 -745
rect 1168 -779 1203 -745
rect 1237 -779 1272 -745
rect 1306 -754 3685 -745
rect 1306 -779 1374 -754
rect -227 -788 1374 -779
rect 1408 -788 1445 -754
rect 1479 -788 1516 -754
rect 1550 -788 1587 -754
rect 1621 -788 1657 -754
rect 1691 -788 1727 -754
rect 1761 -788 1797 -754
rect 1831 -788 1867 -754
rect 1901 -788 1937 -754
rect 1971 -788 2007 -754
rect 2041 -788 2077 -754
rect 2111 -788 2147 -754
rect 2181 -788 2217 -754
rect 2251 -788 2287 -754
rect 2321 -788 2357 -754
rect 2391 -788 2427 -754
rect 2461 -788 2497 -754
rect 2531 -788 2567 -754
rect 2601 -788 2637 -754
rect 2671 -788 2707 -754
rect 2741 -788 2777 -754
rect 2811 -788 2847 -754
rect 2881 -788 2917 -754
rect 2951 -788 2987 -754
rect 3021 -788 3057 -754
rect 3091 -788 3127 -754
rect 3161 -788 3197 -754
rect 3231 -788 3267 -754
rect 3301 -788 3337 -754
rect 3371 -788 3407 -754
rect 3441 -788 3477 -754
rect 3511 -788 3547 -754
rect 3581 -788 3617 -754
rect 3651 -788 3685 -754
rect -227 -817 3685 -788
rect -227 -851 -193 -817
rect -159 -851 -123 -817
rect -89 -851 -53 -817
rect -19 -851 17 -817
rect 51 -851 87 -817
rect 121 -851 157 -817
rect 191 -851 227 -817
rect 261 -851 297 -817
rect 331 -851 367 -817
rect 401 -851 437 -817
rect 471 -851 507 -817
rect 541 -851 577 -817
rect 611 -851 647 -817
rect 681 -851 717 -817
rect 751 -851 787 -817
rect 821 -851 857 -817
rect 891 -851 927 -817
rect 961 -851 996 -817
rect 1030 -851 1065 -817
rect 1099 -851 1134 -817
rect 1168 -851 1203 -817
rect 1237 -851 1272 -817
rect 1306 -824 3685 -817
rect 1306 -851 1374 -824
rect -227 -858 1374 -851
rect 1408 -858 1445 -824
rect 1479 -858 1516 -824
rect 1550 -858 1587 -824
rect 1621 -858 1657 -824
rect 1691 -858 1727 -824
rect 1761 -858 1797 -824
rect 1831 -858 1867 -824
rect 1901 -858 1937 -824
rect 1971 -858 2007 -824
rect 2041 -858 2077 -824
rect 2111 -858 2147 -824
rect 2181 -858 2217 -824
rect 2251 -858 2287 -824
rect 2321 -858 2357 -824
rect 2391 -858 2427 -824
rect 2461 -858 2497 -824
rect 2531 -858 2567 -824
rect 2601 -858 2637 -824
rect 2671 -858 2707 -824
rect 2741 -858 2777 -824
rect 2811 -858 2847 -824
rect 2881 -858 2917 -824
rect 2951 -858 2987 -824
rect 3021 -858 3057 -824
rect 3091 -858 3127 -824
rect 3161 -858 3197 -824
rect 3231 -858 3267 -824
rect 3301 -858 3337 -824
rect 3371 -858 3407 -824
rect 3441 -858 3477 -824
rect 3511 -858 3547 -824
rect 3581 -858 3617 -824
rect 3651 -858 3685 -824
rect -227 -889 3685 -858
rect -227 -923 -193 -889
rect -159 -923 -123 -889
rect -89 -923 -53 -889
rect -19 -923 17 -889
rect 51 -923 87 -889
rect 121 -923 157 -889
rect 191 -923 227 -889
rect 261 -923 297 -889
rect 331 -923 367 -889
rect 401 -923 437 -889
rect 471 -923 507 -889
rect 541 -923 577 -889
rect 611 -923 647 -889
rect 681 -923 717 -889
rect 751 -923 787 -889
rect 821 -923 857 -889
rect 891 -923 927 -889
rect 961 -923 996 -889
rect 1030 -923 1065 -889
rect 1099 -923 1134 -889
rect 1168 -923 1203 -889
rect 1237 -923 1272 -889
rect 1306 -894 3685 -889
rect 1306 -923 1374 -894
rect -227 -928 1374 -923
rect 1408 -928 1445 -894
rect 1479 -928 1516 -894
rect 1550 -928 1587 -894
rect 1621 -928 1657 -894
rect 1691 -928 1727 -894
rect 1761 -928 1797 -894
rect 1831 -928 1867 -894
rect 1901 -928 1937 -894
rect 1971 -928 2007 -894
rect 2041 -928 2077 -894
rect 2111 -928 2147 -894
rect 2181 -928 2217 -894
rect 2251 -928 2287 -894
rect 2321 -928 2357 -894
rect 2391 -928 2427 -894
rect 2461 -928 2497 -894
rect 2531 -928 2567 -894
rect 2601 -928 2637 -894
rect 2671 -928 2707 -894
rect 2741 -928 2777 -894
rect 2811 -928 2847 -894
rect 2881 -928 2917 -894
rect 2951 -928 2987 -894
rect 3021 -928 3057 -894
rect 3091 -928 3127 -894
rect 3161 -928 3197 -894
rect 3231 -928 3267 -894
rect 3301 -928 3337 -894
rect 3371 -928 3407 -894
rect 3441 -928 3477 -894
rect 3511 -928 3547 -894
rect 3581 -928 3617 -894
rect 3651 -928 3685 -894
rect -227 -961 3685 -928
rect -227 -995 -193 -961
rect -159 -995 -123 -961
rect -89 -995 -53 -961
rect -19 -995 17 -961
rect 51 -995 87 -961
rect 121 -995 157 -961
rect 191 -995 227 -961
rect 261 -995 297 -961
rect 331 -995 367 -961
rect 401 -995 437 -961
rect 471 -995 507 -961
rect 541 -995 577 -961
rect 611 -995 647 -961
rect 681 -995 717 -961
rect 751 -995 787 -961
rect 821 -995 857 -961
rect 891 -995 927 -961
rect 961 -995 996 -961
rect 1030 -995 1065 -961
rect 1099 -995 1134 -961
rect 1168 -995 1203 -961
rect 1237 -995 1272 -961
rect 1306 -964 3685 -961
rect 1306 -995 1374 -964
rect -227 -998 1374 -995
rect 1408 -998 1445 -964
rect 1479 -998 1516 -964
rect 1550 -998 1587 -964
rect 1621 -998 1657 -964
rect 1691 -998 1727 -964
rect 1761 -998 1797 -964
rect 1831 -998 1867 -964
rect 1901 -998 1937 -964
rect 1971 -998 2007 -964
rect 2041 -998 2077 -964
rect 2111 -998 2147 -964
rect 2181 -998 2217 -964
rect 2251 -998 2287 -964
rect 2321 -998 2357 -964
rect 2391 -998 2427 -964
rect 2461 -998 2497 -964
rect 2531 -998 2567 -964
rect 2601 -998 2637 -964
rect 2671 -998 2707 -964
rect 2741 -998 2777 -964
rect 2811 -998 2847 -964
rect 2881 -998 2917 -964
rect 2951 -998 2987 -964
rect 3021 -998 3057 -964
rect 3091 -998 3127 -964
rect 3161 -998 3197 -964
rect 3231 -998 3267 -964
rect 3301 -998 3337 -964
rect 3371 -998 3407 -964
rect 3441 -998 3477 -964
rect 3511 -998 3547 -964
rect 3581 -998 3617 -964
rect 3651 -998 3685 -964
rect -227 -1033 3685 -998
rect -227 -1067 -193 -1033
rect -159 -1067 -123 -1033
rect -89 -1067 -53 -1033
rect -19 -1067 17 -1033
rect 51 -1067 87 -1033
rect 121 -1067 157 -1033
rect 191 -1067 227 -1033
rect 261 -1067 297 -1033
rect 331 -1067 367 -1033
rect 401 -1067 437 -1033
rect 471 -1067 507 -1033
rect 541 -1067 577 -1033
rect 611 -1067 647 -1033
rect 681 -1067 717 -1033
rect 751 -1067 787 -1033
rect 821 -1067 857 -1033
rect 891 -1067 927 -1033
rect 961 -1067 996 -1033
rect 1030 -1067 1065 -1033
rect 1099 -1067 1134 -1033
rect 1168 -1067 1203 -1033
rect 1237 -1067 1272 -1033
rect 1306 -1034 3685 -1033
rect 1306 -1067 1374 -1034
rect -227 -1068 1374 -1067
rect 1408 -1068 1445 -1034
rect 1479 -1068 1516 -1034
rect 1550 -1068 1587 -1034
rect 1621 -1068 1657 -1034
rect 1691 -1068 1727 -1034
rect 1761 -1068 1797 -1034
rect 1831 -1068 1867 -1034
rect 1901 -1068 1937 -1034
rect 1971 -1068 2007 -1034
rect 2041 -1068 2077 -1034
rect 2111 -1068 2147 -1034
rect 2181 -1068 2217 -1034
rect 2251 -1068 2287 -1034
rect 2321 -1068 2357 -1034
rect 2391 -1068 2427 -1034
rect 2461 -1068 2497 -1034
rect 2531 -1068 2567 -1034
rect 2601 -1068 2637 -1034
rect 2671 -1068 2707 -1034
rect 2741 -1068 2777 -1034
rect 2811 -1068 2847 -1034
rect 2881 -1068 2917 -1034
rect 2951 -1068 2987 -1034
rect 3021 -1068 3057 -1034
rect 3091 -1068 3127 -1034
rect 3161 -1068 3197 -1034
rect 3231 -1068 3267 -1034
rect 3301 -1068 3337 -1034
rect 3371 -1068 3407 -1034
rect 3441 -1068 3477 -1034
rect 3511 -1068 3547 -1034
rect 3581 -1068 3617 -1034
rect 3651 -1068 3685 -1034
rect -227 -1072 3685 -1068
<< psubdiffcont >>
rect 2596 2171 2630 2205
rect 2669 2171 2703 2205
rect 2741 2171 2775 2205
rect 2813 2171 2847 2205
rect 2885 2171 2919 2205
rect 2957 2171 2991 2205
rect 3029 2171 3063 2205
rect 3101 2171 3135 2205
rect 3173 2171 3207 2205
rect 3245 2171 3279 2205
rect 3317 2171 3351 2205
rect 3389 2171 3423 2205
rect 3461 2171 3495 2205
rect 3533 2171 3567 2205
rect 3605 2171 3639 2205
rect 3677 2171 3711 2205
rect 2596 2103 2630 2137
rect 2669 2103 2703 2137
rect 2741 2103 2775 2137
rect 2813 2103 2847 2137
rect 2885 2103 2919 2137
rect 2957 2103 2991 2137
rect 3029 2103 3063 2137
rect 3101 2103 3135 2137
rect 3173 2103 3207 2137
rect 3245 2103 3279 2137
rect 3317 2103 3351 2137
rect 3389 2103 3423 2137
rect 3461 2103 3495 2137
rect 3533 2103 3567 2137
rect 3605 2103 3639 2137
rect 3677 2103 3711 2137
rect 2596 2035 2630 2069
rect 2669 2035 2703 2069
rect 2741 2035 2775 2069
rect 2813 2035 2847 2069
rect 2885 2035 2919 2069
rect 2957 2035 2991 2069
rect 3029 2035 3063 2069
rect 3101 2035 3135 2069
rect 3173 2035 3207 2069
rect 3245 2035 3279 2069
rect 3317 2035 3351 2069
rect 3389 2035 3423 2069
rect 3461 2035 3495 2069
rect 3533 2035 3567 2069
rect 3605 2035 3639 2069
rect 3677 2035 3711 2069
rect 2596 1967 2630 2001
rect 2669 1967 2703 2001
rect 2741 1967 2775 2001
rect 2813 1967 2847 2001
rect 2885 1967 2919 2001
rect 2957 1967 2991 2001
rect 3029 1967 3063 2001
rect 3101 1967 3135 2001
rect 3173 1967 3207 2001
rect 3245 1967 3279 2001
rect 3317 1967 3351 2001
rect 3389 1967 3423 2001
rect 3461 1967 3495 2001
rect 3533 1967 3567 2001
rect 3605 1967 3639 2001
rect 3677 1967 3711 2001
rect 2579 1899 2613 1933
rect 2648 1899 2682 1933
rect 2717 1899 2751 1933
rect 2786 1899 2820 1933
rect 2855 1899 2889 1933
rect 2924 1899 2958 1933
rect 2993 1899 3027 1933
rect 3062 1899 3096 1933
rect 3131 1899 3165 1933
rect 3200 1899 3234 1933
rect 3269 1899 3303 1933
rect 3338 1899 3372 1933
rect 3407 1899 3441 1933
rect 3476 1899 3510 1933
rect 3545 1899 3579 1933
rect 3613 1899 3647 1933
rect 3681 1899 3715 1933
rect 2579 1819 2613 1853
rect 2648 1819 2682 1853
rect 2717 1819 2751 1853
rect 2786 1819 2820 1853
rect 2855 1819 2889 1853
rect 2924 1819 2958 1853
rect 2993 1819 3027 1853
rect 3062 1819 3096 1853
rect 3131 1819 3165 1853
rect 3200 1819 3234 1853
rect 3269 1819 3303 1853
rect 3338 1819 3372 1853
rect 3407 1819 3441 1853
rect 3476 1819 3510 1853
rect 3545 1819 3579 1853
rect 3613 1819 3647 1853
rect 3681 1819 3715 1853
rect 2579 1739 2613 1773
rect 2648 1739 2682 1773
rect 2717 1739 2751 1773
rect 2786 1739 2820 1773
rect 2855 1739 2889 1773
rect 2924 1739 2958 1773
rect 2993 1739 3027 1773
rect 3062 1739 3096 1773
rect 3131 1739 3165 1773
rect 3200 1739 3234 1773
rect 3269 1739 3303 1773
rect 3338 1739 3372 1773
rect 3407 1739 3441 1773
rect 3476 1739 3510 1773
rect 3545 1739 3579 1773
rect 3613 1739 3647 1773
rect 3681 1739 3715 1773
rect 2579 1659 2613 1693
rect 2648 1659 2682 1693
rect 2717 1659 2751 1693
rect 2786 1659 2820 1693
rect 2855 1659 2889 1693
rect 2924 1659 2958 1693
rect 2993 1659 3027 1693
rect 3062 1659 3096 1693
rect 3131 1659 3165 1693
rect 3200 1659 3234 1693
rect 3269 1659 3303 1693
rect 3338 1659 3372 1693
rect 3407 1659 3441 1693
rect 3476 1659 3510 1693
rect 3545 1659 3579 1693
rect 3613 1659 3647 1693
rect 3681 1659 3715 1693
rect 6102 195 6204 841
rect 6239 195 6341 841
rect 5649 99 5683 133
rect 5934 99 5968 133
rect 6003 99 6037 133
rect 6072 99 6106 133
rect 6141 99 6175 133
rect 6210 99 6244 133
rect 6279 99 6313 133
rect 6348 99 6382 133
rect 6417 99 6451 133
rect 6486 99 6520 133
rect 6555 99 6589 133
rect 6624 99 6658 133
rect 6693 99 6727 133
rect 6762 99 6796 133
rect 6831 99 6865 133
rect 6900 99 6934 133
rect 6969 99 7003 133
rect 7038 99 7072 133
rect 7107 99 7141 133
rect 7176 99 7210 133
rect 7245 99 7279 133
rect 7314 99 7348 133
rect 7383 99 7417 133
rect 7452 99 7486 133
rect 7521 99 7555 133
rect 7590 99 7624 133
rect 7659 99 7693 133
rect 7728 99 7762 133
rect 7797 99 7831 133
rect 7866 99 7900 133
rect 7935 99 7969 133
rect 8004 99 8038 133
rect 8073 99 8107 133
rect 8142 99 8176 133
rect 8211 99 8245 133
rect 8280 99 8314 133
rect 8349 99 8383 133
rect 8418 99 8452 133
rect 8487 99 8521 133
rect 8556 99 8590 133
rect 8625 99 8659 133
rect 8694 99 8728 133
rect 8763 99 8797 133
rect 8832 99 8866 133
rect 8901 99 8935 133
rect 8970 99 9004 133
rect 9039 99 9073 133
rect 9108 99 9142 133
rect 9177 99 9211 133
rect 9246 99 9280 133
rect 9315 99 9349 133
rect 9384 99 9418 133
rect 9453 99 9487 133
rect 9522 99 9556 133
rect 9591 99 9625 133
rect 9660 99 9694 133
rect 9728 99 9762 133
rect 9796 99 9830 133
rect 9864 99 9898 133
rect 9932 99 9966 133
rect 10000 99 10034 133
rect 10068 99 10102 133
rect 10136 99 10170 133
rect 10204 99 10238 133
rect 10272 99 10306 133
rect 10340 99 10374 133
rect 10408 99 10442 133
rect 10476 99 10510 133
rect 10544 99 10578 133
rect 10612 99 10646 133
rect 10680 99 10714 133
rect 10748 99 10782 133
rect 10816 99 10850 133
rect 10884 99 10918 133
rect 10952 99 10986 133
rect 11020 99 11054 133
rect 11088 99 11122 133
rect 11156 99 11190 133
rect 11224 99 11258 133
rect 11292 99 11326 133
rect 11360 99 11394 133
rect 11428 99 11462 133
rect 11496 99 11530 133
rect 11564 99 11598 133
rect 11632 99 11666 133
rect 11700 99 11734 133
rect 11768 99 11802 133
rect 11836 99 11870 133
rect 11904 99 11938 133
rect 11972 99 12006 133
rect 12040 99 12074 133
rect 1374 -158 1408 -124
rect 1445 -158 1479 -124
rect 1516 -158 1550 -124
rect 1587 -158 1621 -124
rect 1657 -158 1691 -124
rect 1727 -158 1761 -124
rect 1797 -158 1831 -124
rect 1867 -158 1901 -124
rect 1937 -158 1971 -124
rect 2007 -158 2041 -124
rect 2077 -158 2111 -124
rect 2147 -158 2181 -124
rect 2217 -158 2251 -124
rect 2287 -158 2321 -124
rect 2357 -158 2391 -124
rect 2427 -158 2461 -124
rect 2497 -158 2531 -124
rect 2567 -158 2601 -124
rect 2637 -158 2671 -124
rect 2707 -158 2741 -124
rect 2777 -158 2811 -124
rect 2847 -158 2881 -124
rect 2917 -158 2951 -124
rect 2987 -158 3021 -124
rect 3057 -158 3091 -124
rect 3127 -158 3161 -124
rect 3197 -158 3231 -124
rect 3267 -158 3301 -124
rect 3337 -158 3371 -124
rect 3407 -158 3441 -124
rect 3477 -158 3511 -124
rect 3547 -158 3581 -124
rect 3617 -158 3651 -124
rect 1374 -228 1408 -194
rect 1445 -228 1479 -194
rect 1516 -228 1550 -194
rect 1587 -228 1621 -194
rect 1657 -228 1691 -194
rect 1727 -228 1761 -194
rect 1797 -228 1831 -194
rect 1867 -228 1901 -194
rect 1937 -228 1971 -194
rect 2007 -228 2041 -194
rect 2077 -228 2111 -194
rect 2147 -228 2181 -194
rect 2217 -228 2251 -194
rect 2287 -228 2321 -194
rect 2357 -228 2391 -194
rect 2427 -228 2461 -194
rect 2497 -228 2531 -194
rect 2567 -228 2601 -194
rect 2637 -228 2671 -194
rect 2707 -228 2741 -194
rect 2777 -228 2811 -194
rect 2847 -228 2881 -194
rect 2917 -228 2951 -194
rect 2987 -228 3021 -194
rect 3057 -228 3091 -194
rect 3127 -228 3161 -194
rect 3197 -228 3231 -194
rect 3267 -228 3301 -194
rect 3337 -228 3371 -194
rect 3407 -228 3441 -194
rect 3477 -228 3511 -194
rect 3547 -228 3581 -194
rect 3617 -228 3651 -194
rect 1374 -298 1408 -264
rect 1445 -298 1479 -264
rect 1516 -298 1550 -264
rect 1587 -298 1621 -264
rect 1657 -298 1691 -264
rect 1727 -298 1761 -264
rect 1797 -298 1831 -264
rect 1867 -298 1901 -264
rect 1937 -298 1971 -264
rect 2007 -298 2041 -264
rect 2077 -298 2111 -264
rect 2147 -298 2181 -264
rect 2217 -298 2251 -264
rect 2287 -298 2321 -264
rect 2357 -298 2391 -264
rect 2427 -298 2461 -264
rect 2497 -298 2531 -264
rect 2567 -298 2601 -264
rect 2637 -298 2671 -264
rect 2707 -298 2741 -264
rect 2777 -298 2811 -264
rect 2847 -298 2881 -264
rect 2917 -298 2951 -264
rect 2987 -298 3021 -264
rect 3057 -298 3091 -264
rect 3127 -298 3161 -264
rect 3197 -298 3231 -264
rect 3267 -298 3301 -264
rect 3337 -298 3371 -264
rect 3407 -298 3441 -264
rect 3477 -298 3511 -264
rect 3547 -298 3581 -264
rect 3617 -298 3651 -264
rect -193 -347 -159 -313
rect -123 -347 -89 -313
rect -53 -347 -19 -313
rect 17 -347 51 -313
rect 87 -347 121 -313
rect 157 -347 191 -313
rect 227 -347 261 -313
rect 297 -347 331 -313
rect 367 -347 401 -313
rect 437 -347 471 -313
rect 507 -347 541 -313
rect 577 -347 611 -313
rect 647 -347 681 -313
rect 717 -347 751 -313
rect 787 -347 821 -313
rect 857 -347 891 -313
rect 927 -347 961 -313
rect 996 -347 1030 -313
rect 1065 -347 1099 -313
rect 1134 -347 1168 -313
rect 1203 -347 1237 -313
rect 1272 -347 1306 -313
rect 1374 -368 1408 -334
rect 1445 -368 1479 -334
rect 1516 -368 1550 -334
rect 1587 -368 1621 -334
rect 1657 -368 1691 -334
rect 1727 -368 1761 -334
rect 1797 -368 1831 -334
rect 1867 -368 1901 -334
rect 1937 -368 1971 -334
rect 2007 -368 2041 -334
rect 2077 -368 2111 -334
rect 2147 -368 2181 -334
rect 2217 -368 2251 -334
rect 2287 -368 2321 -334
rect 2357 -368 2391 -334
rect 2427 -368 2461 -334
rect 2497 -368 2531 -334
rect 2567 -368 2601 -334
rect 2637 -368 2671 -334
rect 2707 -368 2741 -334
rect 2777 -368 2811 -334
rect 2847 -368 2881 -334
rect 2917 -368 2951 -334
rect 2987 -368 3021 -334
rect 3057 -368 3091 -334
rect 3127 -368 3161 -334
rect 3197 -368 3231 -334
rect 3267 -368 3301 -334
rect 3337 -368 3371 -334
rect 3407 -368 3441 -334
rect 3477 -368 3511 -334
rect 3547 -368 3581 -334
rect 3617 -368 3651 -334
rect -193 -419 -159 -385
rect -123 -419 -89 -385
rect -53 -419 -19 -385
rect 17 -419 51 -385
rect 87 -419 121 -385
rect 157 -419 191 -385
rect 227 -419 261 -385
rect 297 -419 331 -385
rect 367 -419 401 -385
rect 437 -419 471 -385
rect 507 -419 541 -385
rect 577 -419 611 -385
rect 647 -419 681 -385
rect 717 -419 751 -385
rect 787 -419 821 -385
rect 857 -419 891 -385
rect 927 -419 961 -385
rect 996 -419 1030 -385
rect 1065 -419 1099 -385
rect 1134 -419 1168 -385
rect 1203 -419 1237 -385
rect 1272 -419 1306 -385
rect 1374 -438 1408 -404
rect 1445 -438 1479 -404
rect 1516 -438 1550 -404
rect 1587 -438 1621 -404
rect 1657 -438 1691 -404
rect 1727 -438 1761 -404
rect 1797 -438 1831 -404
rect 1867 -438 1901 -404
rect 1937 -438 1971 -404
rect 2007 -438 2041 -404
rect 2077 -438 2111 -404
rect 2147 -438 2181 -404
rect 2217 -438 2251 -404
rect 2287 -438 2321 -404
rect 2357 -438 2391 -404
rect 2427 -438 2461 -404
rect 2497 -438 2531 -404
rect 2567 -438 2601 -404
rect 2637 -438 2671 -404
rect 2707 -438 2741 -404
rect 2777 -438 2811 -404
rect 2847 -438 2881 -404
rect 2917 -438 2951 -404
rect 2987 -438 3021 -404
rect 3057 -438 3091 -404
rect 3127 -438 3161 -404
rect 3197 -438 3231 -404
rect 3267 -438 3301 -404
rect 3337 -438 3371 -404
rect 3407 -438 3441 -404
rect 3477 -438 3511 -404
rect 3547 -438 3581 -404
rect 3617 -438 3651 -404
rect -193 -491 -159 -457
rect -123 -491 -89 -457
rect -53 -491 -19 -457
rect 17 -491 51 -457
rect 87 -491 121 -457
rect 157 -491 191 -457
rect 227 -491 261 -457
rect 297 -491 331 -457
rect 367 -491 401 -457
rect 437 -491 471 -457
rect 507 -491 541 -457
rect 577 -491 611 -457
rect 647 -491 681 -457
rect 717 -491 751 -457
rect 787 -491 821 -457
rect 857 -491 891 -457
rect 927 -491 961 -457
rect 996 -491 1030 -457
rect 1065 -491 1099 -457
rect 1134 -491 1168 -457
rect 1203 -491 1237 -457
rect 1272 -491 1306 -457
rect 1374 -508 1408 -474
rect 1445 -508 1479 -474
rect 1516 -508 1550 -474
rect 1587 -508 1621 -474
rect 1657 -508 1691 -474
rect 1727 -508 1761 -474
rect 1797 -508 1831 -474
rect 1867 -508 1901 -474
rect 1937 -508 1971 -474
rect 2007 -508 2041 -474
rect 2077 -508 2111 -474
rect 2147 -508 2181 -474
rect 2217 -508 2251 -474
rect 2287 -508 2321 -474
rect 2357 -508 2391 -474
rect 2427 -508 2461 -474
rect 2497 -508 2531 -474
rect 2567 -508 2601 -474
rect 2637 -508 2671 -474
rect 2707 -508 2741 -474
rect 2777 -508 2811 -474
rect 2847 -508 2881 -474
rect 2917 -508 2951 -474
rect 2987 -508 3021 -474
rect 3057 -508 3091 -474
rect 3127 -508 3161 -474
rect 3197 -508 3231 -474
rect 3267 -508 3301 -474
rect 3337 -508 3371 -474
rect 3407 -508 3441 -474
rect 3477 -508 3511 -474
rect 3547 -508 3581 -474
rect 3617 -508 3651 -474
rect -193 -563 -159 -529
rect -123 -563 -89 -529
rect -53 -563 -19 -529
rect 17 -563 51 -529
rect 87 -563 121 -529
rect 157 -563 191 -529
rect 227 -563 261 -529
rect 297 -563 331 -529
rect 367 -563 401 -529
rect 437 -563 471 -529
rect 507 -563 541 -529
rect 577 -563 611 -529
rect 647 -563 681 -529
rect 717 -563 751 -529
rect 787 -563 821 -529
rect 857 -563 891 -529
rect 927 -563 961 -529
rect 996 -563 1030 -529
rect 1065 -563 1099 -529
rect 1134 -563 1168 -529
rect 1203 -563 1237 -529
rect 1272 -563 1306 -529
rect 1374 -578 1408 -544
rect 1445 -578 1479 -544
rect 1516 -578 1550 -544
rect 1587 -578 1621 -544
rect 1657 -578 1691 -544
rect 1727 -578 1761 -544
rect 1797 -578 1831 -544
rect 1867 -578 1901 -544
rect 1937 -578 1971 -544
rect 2007 -578 2041 -544
rect 2077 -578 2111 -544
rect 2147 -578 2181 -544
rect 2217 -578 2251 -544
rect 2287 -578 2321 -544
rect 2357 -578 2391 -544
rect 2427 -578 2461 -544
rect 2497 -578 2531 -544
rect 2567 -578 2601 -544
rect 2637 -578 2671 -544
rect 2707 -578 2741 -544
rect 2777 -578 2811 -544
rect 2847 -578 2881 -544
rect 2917 -578 2951 -544
rect 2987 -578 3021 -544
rect 3057 -578 3091 -544
rect 3127 -578 3161 -544
rect 3197 -578 3231 -544
rect 3267 -578 3301 -544
rect 3337 -578 3371 -544
rect 3407 -578 3441 -544
rect 3477 -578 3511 -544
rect 3547 -578 3581 -544
rect 3617 -578 3651 -544
rect -193 -635 -159 -601
rect -123 -635 -89 -601
rect -53 -635 -19 -601
rect 17 -635 51 -601
rect 87 -635 121 -601
rect 157 -635 191 -601
rect 227 -635 261 -601
rect 297 -635 331 -601
rect 367 -635 401 -601
rect 437 -635 471 -601
rect 507 -635 541 -601
rect 577 -635 611 -601
rect 647 -635 681 -601
rect 717 -635 751 -601
rect 787 -635 821 -601
rect 857 -635 891 -601
rect 927 -635 961 -601
rect 996 -635 1030 -601
rect 1065 -635 1099 -601
rect 1134 -635 1168 -601
rect 1203 -635 1237 -601
rect 1272 -635 1306 -601
rect 1374 -648 1408 -614
rect 1445 -648 1479 -614
rect 1516 -648 1550 -614
rect 1587 -648 1621 -614
rect 1657 -648 1691 -614
rect 1727 -648 1761 -614
rect 1797 -648 1831 -614
rect 1867 -648 1901 -614
rect 1937 -648 1971 -614
rect 2007 -648 2041 -614
rect 2077 -648 2111 -614
rect 2147 -648 2181 -614
rect 2217 -648 2251 -614
rect 2287 -648 2321 -614
rect 2357 -648 2391 -614
rect 2427 -648 2461 -614
rect 2497 -648 2531 -614
rect 2567 -648 2601 -614
rect 2637 -648 2671 -614
rect 2707 -648 2741 -614
rect 2777 -648 2811 -614
rect 2847 -648 2881 -614
rect 2917 -648 2951 -614
rect 2987 -648 3021 -614
rect 3057 -648 3091 -614
rect 3127 -648 3161 -614
rect 3197 -648 3231 -614
rect 3267 -648 3301 -614
rect 3337 -648 3371 -614
rect 3407 -648 3441 -614
rect 3477 -648 3511 -614
rect 3547 -648 3581 -614
rect 3617 -648 3651 -614
rect -193 -707 -159 -673
rect -123 -707 -89 -673
rect -53 -707 -19 -673
rect 17 -707 51 -673
rect 87 -707 121 -673
rect 157 -707 191 -673
rect 227 -707 261 -673
rect 297 -707 331 -673
rect 367 -707 401 -673
rect 437 -707 471 -673
rect 507 -707 541 -673
rect 577 -707 611 -673
rect 647 -707 681 -673
rect 717 -707 751 -673
rect 787 -707 821 -673
rect 857 -707 891 -673
rect 927 -707 961 -673
rect 996 -707 1030 -673
rect 1065 -707 1099 -673
rect 1134 -707 1168 -673
rect 1203 -707 1237 -673
rect 1272 -707 1306 -673
rect 1374 -718 1408 -684
rect 1445 -718 1479 -684
rect 1516 -718 1550 -684
rect 1587 -718 1621 -684
rect 1657 -718 1691 -684
rect 1727 -718 1761 -684
rect 1797 -718 1831 -684
rect 1867 -718 1901 -684
rect 1937 -718 1971 -684
rect 2007 -718 2041 -684
rect 2077 -718 2111 -684
rect 2147 -718 2181 -684
rect 2217 -718 2251 -684
rect 2287 -718 2321 -684
rect 2357 -718 2391 -684
rect 2427 -718 2461 -684
rect 2497 -718 2531 -684
rect 2567 -718 2601 -684
rect 2637 -718 2671 -684
rect 2707 -718 2741 -684
rect 2777 -718 2811 -684
rect 2847 -718 2881 -684
rect 2917 -718 2951 -684
rect 2987 -718 3021 -684
rect 3057 -718 3091 -684
rect 3127 -718 3161 -684
rect 3197 -718 3231 -684
rect 3267 -718 3301 -684
rect 3337 -718 3371 -684
rect 3407 -718 3441 -684
rect 3477 -718 3511 -684
rect 3547 -718 3581 -684
rect 3617 -718 3651 -684
rect -193 -779 -159 -745
rect -123 -779 -89 -745
rect -53 -779 -19 -745
rect 17 -779 51 -745
rect 87 -779 121 -745
rect 157 -779 191 -745
rect 227 -779 261 -745
rect 297 -779 331 -745
rect 367 -779 401 -745
rect 437 -779 471 -745
rect 507 -779 541 -745
rect 577 -779 611 -745
rect 647 -779 681 -745
rect 717 -779 751 -745
rect 787 -779 821 -745
rect 857 -779 891 -745
rect 927 -779 961 -745
rect 996 -779 1030 -745
rect 1065 -779 1099 -745
rect 1134 -779 1168 -745
rect 1203 -779 1237 -745
rect 1272 -779 1306 -745
rect 1374 -788 1408 -754
rect 1445 -788 1479 -754
rect 1516 -788 1550 -754
rect 1587 -788 1621 -754
rect 1657 -788 1691 -754
rect 1727 -788 1761 -754
rect 1797 -788 1831 -754
rect 1867 -788 1901 -754
rect 1937 -788 1971 -754
rect 2007 -788 2041 -754
rect 2077 -788 2111 -754
rect 2147 -788 2181 -754
rect 2217 -788 2251 -754
rect 2287 -788 2321 -754
rect 2357 -788 2391 -754
rect 2427 -788 2461 -754
rect 2497 -788 2531 -754
rect 2567 -788 2601 -754
rect 2637 -788 2671 -754
rect 2707 -788 2741 -754
rect 2777 -788 2811 -754
rect 2847 -788 2881 -754
rect 2917 -788 2951 -754
rect 2987 -788 3021 -754
rect 3057 -788 3091 -754
rect 3127 -788 3161 -754
rect 3197 -788 3231 -754
rect 3267 -788 3301 -754
rect 3337 -788 3371 -754
rect 3407 -788 3441 -754
rect 3477 -788 3511 -754
rect 3547 -788 3581 -754
rect 3617 -788 3651 -754
rect -193 -851 -159 -817
rect -123 -851 -89 -817
rect -53 -851 -19 -817
rect 17 -851 51 -817
rect 87 -851 121 -817
rect 157 -851 191 -817
rect 227 -851 261 -817
rect 297 -851 331 -817
rect 367 -851 401 -817
rect 437 -851 471 -817
rect 507 -851 541 -817
rect 577 -851 611 -817
rect 647 -851 681 -817
rect 717 -851 751 -817
rect 787 -851 821 -817
rect 857 -851 891 -817
rect 927 -851 961 -817
rect 996 -851 1030 -817
rect 1065 -851 1099 -817
rect 1134 -851 1168 -817
rect 1203 -851 1237 -817
rect 1272 -851 1306 -817
rect 1374 -858 1408 -824
rect 1445 -858 1479 -824
rect 1516 -858 1550 -824
rect 1587 -858 1621 -824
rect 1657 -858 1691 -824
rect 1727 -858 1761 -824
rect 1797 -858 1831 -824
rect 1867 -858 1901 -824
rect 1937 -858 1971 -824
rect 2007 -858 2041 -824
rect 2077 -858 2111 -824
rect 2147 -858 2181 -824
rect 2217 -858 2251 -824
rect 2287 -858 2321 -824
rect 2357 -858 2391 -824
rect 2427 -858 2461 -824
rect 2497 -858 2531 -824
rect 2567 -858 2601 -824
rect 2637 -858 2671 -824
rect 2707 -858 2741 -824
rect 2777 -858 2811 -824
rect 2847 -858 2881 -824
rect 2917 -858 2951 -824
rect 2987 -858 3021 -824
rect 3057 -858 3091 -824
rect 3127 -858 3161 -824
rect 3197 -858 3231 -824
rect 3267 -858 3301 -824
rect 3337 -858 3371 -824
rect 3407 -858 3441 -824
rect 3477 -858 3511 -824
rect 3547 -858 3581 -824
rect 3617 -858 3651 -824
rect -193 -923 -159 -889
rect -123 -923 -89 -889
rect -53 -923 -19 -889
rect 17 -923 51 -889
rect 87 -923 121 -889
rect 157 -923 191 -889
rect 227 -923 261 -889
rect 297 -923 331 -889
rect 367 -923 401 -889
rect 437 -923 471 -889
rect 507 -923 541 -889
rect 577 -923 611 -889
rect 647 -923 681 -889
rect 717 -923 751 -889
rect 787 -923 821 -889
rect 857 -923 891 -889
rect 927 -923 961 -889
rect 996 -923 1030 -889
rect 1065 -923 1099 -889
rect 1134 -923 1168 -889
rect 1203 -923 1237 -889
rect 1272 -923 1306 -889
rect 1374 -928 1408 -894
rect 1445 -928 1479 -894
rect 1516 -928 1550 -894
rect 1587 -928 1621 -894
rect 1657 -928 1691 -894
rect 1727 -928 1761 -894
rect 1797 -928 1831 -894
rect 1867 -928 1901 -894
rect 1937 -928 1971 -894
rect 2007 -928 2041 -894
rect 2077 -928 2111 -894
rect 2147 -928 2181 -894
rect 2217 -928 2251 -894
rect 2287 -928 2321 -894
rect 2357 -928 2391 -894
rect 2427 -928 2461 -894
rect 2497 -928 2531 -894
rect 2567 -928 2601 -894
rect 2637 -928 2671 -894
rect 2707 -928 2741 -894
rect 2777 -928 2811 -894
rect 2847 -928 2881 -894
rect 2917 -928 2951 -894
rect 2987 -928 3021 -894
rect 3057 -928 3091 -894
rect 3127 -928 3161 -894
rect 3197 -928 3231 -894
rect 3267 -928 3301 -894
rect 3337 -928 3371 -894
rect 3407 -928 3441 -894
rect 3477 -928 3511 -894
rect 3547 -928 3581 -894
rect 3617 -928 3651 -894
rect -193 -995 -159 -961
rect -123 -995 -89 -961
rect -53 -995 -19 -961
rect 17 -995 51 -961
rect 87 -995 121 -961
rect 157 -995 191 -961
rect 227 -995 261 -961
rect 297 -995 331 -961
rect 367 -995 401 -961
rect 437 -995 471 -961
rect 507 -995 541 -961
rect 577 -995 611 -961
rect 647 -995 681 -961
rect 717 -995 751 -961
rect 787 -995 821 -961
rect 857 -995 891 -961
rect 927 -995 961 -961
rect 996 -995 1030 -961
rect 1065 -995 1099 -961
rect 1134 -995 1168 -961
rect 1203 -995 1237 -961
rect 1272 -995 1306 -961
rect 1374 -998 1408 -964
rect 1445 -998 1479 -964
rect 1516 -998 1550 -964
rect 1587 -998 1621 -964
rect 1657 -998 1691 -964
rect 1727 -998 1761 -964
rect 1797 -998 1831 -964
rect 1867 -998 1901 -964
rect 1937 -998 1971 -964
rect 2007 -998 2041 -964
rect 2077 -998 2111 -964
rect 2147 -998 2181 -964
rect 2217 -998 2251 -964
rect 2287 -998 2321 -964
rect 2357 -998 2391 -964
rect 2427 -998 2461 -964
rect 2497 -998 2531 -964
rect 2567 -998 2601 -964
rect 2637 -998 2671 -964
rect 2707 -998 2741 -964
rect 2777 -998 2811 -964
rect 2847 -998 2881 -964
rect 2917 -998 2951 -964
rect 2987 -998 3021 -964
rect 3057 -998 3091 -964
rect 3127 -998 3161 -964
rect 3197 -998 3231 -964
rect 3267 -998 3301 -964
rect 3337 -998 3371 -964
rect 3407 -998 3441 -964
rect 3477 -998 3511 -964
rect 3547 -998 3581 -964
rect 3617 -998 3651 -964
rect -193 -1067 -159 -1033
rect -123 -1067 -89 -1033
rect -53 -1067 -19 -1033
rect 17 -1067 51 -1033
rect 87 -1067 121 -1033
rect 157 -1067 191 -1033
rect 227 -1067 261 -1033
rect 297 -1067 331 -1033
rect 367 -1067 401 -1033
rect 437 -1067 471 -1033
rect 507 -1067 541 -1033
rect 577 -1067 611 -1033
rect 647 -1067 681 -1033
rect 717 -1067 751 -1033
rect 787 -1067 821 -1033
rect 857 -1067 891 -1033
rect 927 -1067 961 -1033
rect 996 -1067 1030 -1033
rect 1065 -1067 1099 -1033
rect 1134 -1067 1168 -1033
rect 1203 -1067 1237 -1033
rect 1272 -1067 1306 -1033
rect 1374 -1068 1408 -1034
rect 1445 -1068 1479 -1034
rect 1516 -1068 1550 -1034
rect 1587 -1068 1621 -1034
rect 1657 -1068 1691 -1034
rect 1727 -1068 1761 -1034
rect 1797 -1068 1831 -1034
rect 1867 -1068 1901 -1034
rect 1937 -1068 1971 -1034
rect 2007 -1068 2041 -1034
rect 2077 -1068 2111 -1034
rect 2147 -1068 2181 -1034
rect 2217 -1068 2251 -1034
rect 2287 -1068 2321 -1034
rect 2357 -1068 2391 -1034
rect 2427 -1068 2461 -1034
rect 2497 -1068 2531 -1034
rect 2567 -1068 2601 -1034
rect 2637 -1068 2671 -1034
rect 2707 -1068 2741 -1034
rect 2777 -1068 2811 -1034
rect 2847 -1068 2881 -1034
rect 2917 -1068 2951 -1034
rect 2987 -1068 3021 -1034
rect 3057 -1068 3091 -1034
rect 3127 -1068 3161 -1034
rect 3197 -1068 3231 -1034
rect 3267 -1068 3301 -1034
rect 3337 -1068 3371 -1034
rect 3407 -1068 3441 -1034
rect 3477 -1068 3511 -1034
rect 3547 -1068 3581 -1034
rect 3617 -1068 3651 -1034
<< poly >>
rect 28 1866 128 1881
rect 28 1850 228 1866
rect 28 1816 178 1850
rect 212 1816 228 1850
rect 28 1782 228 1816
rect 28 1762 178 1782
rect 162 1748 178 1762
rect 212 1748 228 1782
rect 162 1732 228 1748
<< polycont >>
rect 178 1816 212 1850
rect 178 1748 212 1782
<< locali >>
rect 2537 2171 2596 2205
rect 2630 2171 2669 2205
rect 2703 2171 2741 2205
rect 2775 2171 2813 2205
rect 2847 2171 2885 2205
rect 2919 2171 2957 2205
rect 2991 2171 3029 2205
rect 3063 2171 3101 2205
rect 3135 2171 3173 2205
rect 3207 2171 3245 2205
rect 3279 2171 3317 2205
rect 3351 2171 3389 2205
rect 3423 2171 3461 2205
rect 3495 2171 3533 2205
rect 3567 2171 3605 2205
rect 3639 2171 3677 2205
rect 3711 2171 3759 2205
rect 139 1850 214 1866
rect 139 1816 178 1850
rect 212 1816 214 1850
rect 139 1782 214 1816
rect 139 1748 178 1782
rect 212 1748 214 1782
rect 139 1482 214 1748
rect 493 1583 588 2145
rect 2537 2137 3759 2171
rect 2537 2103 2596 2137
rect 2630 2103 2669 2137
rect 2703 2103 2741 2137
rect 2775 2103 2813 2137
rect 2847 2103 2885 2137
rect 2919 2103 2957 2137
rect 2991 2103 3029 2137
rect 3063 2103 3101 2137
rect 3135 2103 3173 2137
rect 3207 2103 3245 2137
rect 3279 2103 3317 2137
rect 3351 2103 3389 2137
rect 3423 2103 3461 2137
rect 3495 2103 3533 2137
rect 3567 2103 3605 2137
rect 3639 2103 3677 2137
rect 3711 2103 3759 2137
rect 2537 2069 3759 2103
rect 2537 2035 2596 2069
rect 2630 2035 2669 2069
rect 2703 2035 2741 2069
rect 2775 2035 2813 2069
rect 2847 2035 2885 2069
rect 2919 2035 2957 2069
rect 2991 2035 3029 2069
rect 3063 2035 3101 2069
rect 3135 2035 3173 2069
rect 3207 2035 3245 2069
rect 3279 2035 3317 2069
rect 3351 2035 3389 2069
rect 3423 2035 3461 2069
rect 3495 2035 3533 2069
rect 3567 2035 3605 2069
rect 3639 2035 3677 2069
rect 3711 2035 3759 2069
rect 2537 2001 3759 2035
rect 2537 1999 2596 2001
rect 2630 1999 2669 2001
rect 2703 1999 2741 2001
rect 2775 1999 2813 2001
rect 2847 1999 2885 2001
rect 2919 1999 2957 2001
rect 2991 1999 3029 2001
rect 3063 1999 3101 2001
rect 3135 1999 3173 2001
rect 3207 1999 3245 2001
rect 3279 1999 3317 2001
rect 3351 1999 3389 2001
rect 3423 1999 3461 2001
rect 3495 1999 3533 2001
rect 3567 1999 3605 2001
rect 3639 1999 3677 2001
rect 2537 1965 2582 1999
rect 2630 1967 2655 1999
rect 2703 1967 2728 1999
rect 2775 1967 2801 1999
rect 2847 1967 2874 1999
rect 2919 1967 2947 1999
rect 2991 1967 3020 1999
rect 3063 1967 3092 1999
rect 3135 1967 3164 1999
rect 3207 1967 3236 1999
rect 3279 1967 3308 1999
rect 3351 1967 3380 1999
rect 3423 1967 3452 1999
rect 3495 1967 3524 1999
rect 3567 1967 3596 1999
rect 3639 1967 3668 1999
rect 3711 1967 3759 2001
rect 2616 1965 2655 1967
rect 2689 1965 2728 1967
rect 2762 1965 2801 1967
rect 2835 1965 2874 1967
rect 2908 1965 2947 1967
rect 2981 1965 3020 1967
rect 3054 1965 3092 1967
rect 3126 1965 3164 1967
rect 3198 1965 3236 1967
rect 3270 1965 3308 1967
rect 3342 1965 3380 1967
rect 3414 1965 3452 1967
rect 3486 1965 3524 1967
rect 3558 1965 3596 1967
rect 3630 1965 3668 1967
rect 3702 1965 3759 1967
rect 2537 1933 3759 1965
rect 2537 1899 2579 1933
rect 2613 1915 2648 1933
rect 2682 1915 2717 1933
rect 2751 1915 2786 1933
rect 2820 1915 2855 1933
rect 2889 1915 2924 1933
rect 2958 1915 2993 1933
rect 3027 1915 3062 1933
rect 3096 1915 3131 1933
rect 3165 1915 3200 1933
rect 2616 1899 2648 1915
rect 2689 1899 2717 1915
rect 2762 1899 2786 1915
rect 2835 1899 2855 1915
rect 2908 1899 2924 1915
rect 2981 1899 2993 1915
rect 3054 1899 3062 1915
rect 3126 1899 3131 1915
rect 3198 1899 3200 1915
rect 3234 1915 3269 1933
rect 3303 1915 3338 1933
rect 3372 1915 3407 1933
rect 3441 1915 3476 1933
rect 3510 1915 3545 1933
rect 3579 1915 3613 1933
rect 3647 1915 3681 1933
rect 3234 1899 3236 1915
rect 3303 1899 3308 1915
rect 3372 1899 3380 1915
rect 3441 1899 3452 1915
rect 3510 1899 3524 1915
rect 3579 1899 3596 1915
rect 3647 1899 3668 1915
rect 3715 1899 3759 1933
rect 2537 1881 2582 1899
rect 2616 1881 2655 1899
rect 2689 1881 2728 1899
rect 2762 1881 2801 1899
rect 2835 1881 2874 1899
rect 2908 1881 2947 1899
rect 2981 1881 3020 1899
rect 3054 1881 3092 1899
rect 3126 1881 3164 1899
rect 3198 1881 3236 1899
rect 3270 1881 3308 1899
rect 3342 1881 3380 1899
rect 3414 1881 3452 1899
rect 3486 1881 3524 1899
rect 3558 1881 3596 1899
rect 3630 1881 3668 1899
rect 3702 1881 3759 1899
rect 2537 1853 3759 1881
rect 2537 1819 2579 1853
rect 2613 1819 2648 1853
rect 2682 1819 2717 1853
rect 2751 1819 2786 1853
rect 2820 1819 2855 1853
rect 2889 1819 2924 1853
rect 2958 1819 2993 1853
rect 3027 1819 3062 1853
rect 3096 1819 3131 1853
rect 3165 1819 3200 1853
rect 3234 1819 3269 1853
rect 3303 1819 3338 1853
rect 3372 1819 3407 1853
rect 3441 1819 3476 1853
rect 3510 1819 3545 1853
rect 3579 1819 3613 1853
rect 3647 1819 3681 1853
rect 3715 1819 3759 1853
rect 2537 1773 3759 1819
rect 2537 1739 2579 1773
rect 2613 1739 2648 1773
rect 2682 1739 2717 1773
rect 2751 1739 2786 1773
rect 2820 1739 2855 1773
rect 2889 1739 2924 1773
rect 2958 1739 2993 1773
rect 3027 1739 3062 1773
rect 3096 1739 3131 1773
rect 3165 1739 3200 1773
rect 3234 1739 3269 1773
rect 3303 1739 3338 1773
rect 3372 1739 3407 1773
rect 3441 1739 3476 1773
rect 3510 1739 3545 1773
rect 3579 1739 3613 1773
rect 3647 1739 3681 1773
rect 3715 1739 3759 1773
rect 2537 1693 3759 1739
rect 2537 1659 2579 1693
rect 2613 1659 2648 1693
rect 2682 1659 2717 1693
rect 2751 1659 2786 1693
rect 2820 1659 2855 1693
rect 2889 1659 2924 1693
rect 2958 1659 2993 1693
rect 3027 1659 3062 1693
rect 3096 1659 3131 1693
rect 3165 1659 3200 1693
rect 3234 1659 3269 1693
rect 3303 1659 3338 1693
rect 3372 1659 3407 1693
rect 3441 1659 3476 1693
rect 3510 1659 3545 1693
rect 3579 1659 3613 1693
rect 3647 1659 3681 1693
rect 3715 1659 3759 1693
rect 2537 1625 3759 1659
rect 522 1549 560 1583
rect 413 1188 448 1234
rect 5831 1167 5869 1201
rect 849 1052 923 1086
rect 849 1018 868 1052
rect 902 1018 923 1052
rect 849 980 923 1018
rect 849 946 868 980
rect 902 946 923 980
rect 849 267 923 946
rect 5197 624 5271 1086
rect 5197 590 5218 624
rect 5252 590 5271 624
rect 5197 552 5271 590
rect 5197 518 5218 552
rect 5252 518 5271 552
rect 5197 267 5271 518
rect 5373 1040 5447 1086
rect 5373 1006 5394 1040
rect 5428 1006 5447 1040
rect 5373 968 5447 1006
rect 7050 1002 7084 1040
rect 5373 934 5394 968
rect 5428 934 5447 968
rect 5373 267 5447 934
rect 6009 841 6375 862
rect 6009 315 6102 841
rect 6069 195 6102 315
rect 6204 195 6239 841
rect 6341 195 6375 841
rect 6690 205 6724 275
rect 7152 205 7186 275
rect 7504 205 7538 275
rect 7856 205 7890 275
rect 8780 205 8814 275
rect 9132 205 9166 275
rect 9484 205 9518 275
rect 9836 205 9870 275
rect 10188 205 10222 275
rect 10540 205 10574 275
rect 10892 205 10926 275
rect 11244 205 11278 275
rect 11596 205 11630 275
rect 11948 205 11982 275
rect 6069 175 6375 195
rect 6069 133 12098 175
rect 5565 99 5620 133
rect 5625 99 5649 133
rect 5683 99 5934 133
rect 5968 99 6003 133
rect 6037 99 6072 133
rect 6106 99 6141 133
rect 6175 99 6210 133
rect 6244 99 6279 133
rect 6313 99 6348 133
rect 6382 99 6417 133
rect 6451 99 6486 133
rect 6520 99 6555 133
rect 6589 99 6624 133
rect 6658 99 6693 133
rect 6727 99 6762 133
rect 6796 99 6831 133
rect 6865 99 6900 133
rect 6934 99 6969 133
rect 7003 99 7038 133
rect 7072 99 7107 133
rect 7141 99 7176 133
rect 7210 99 7245 133
rect 7279 99 7314 133
rect 7348 99 7383 133
rect 7417 99 7452 133
rect 7486 99 7521 133
rect 7555 99 7590 133
rect 7624 99 7659 133
rect 7693 99 7728 133
rect 7762 99 7797 133
rect 7831 99 7866 133
rect 7900 99 7935 133
rect 7969 99 8004 133
rect 8038 99 8073 133
rect 8107 99 8142 133
rect 8176 99 8211 133
rect 8245 99 8280 133
rect 8314 99 8349 133
rect 8383 99 8418 133
rect 8452 99 8487 133
rect 8521 99 8556 133
rect 8590 99 8625 133
rect 8659 99 8694 133
rect 8728 99 8763 133
rect 8797 99 8832 133
rect 8866 99 8901 133
rect 8935 99 8970 133
rect 9004 99 9039 133
rect 9073 99 9108 133
rect 9142 99 9177 133
rect 9211 99 9246 133
rect 9280 99 9315 133
rect 9349 99 9384 133
rect 9418 99 9453 133
rect 9487 99 9522 133
rect 9556 99 9591 133
rect 9625 99 9660 133
rect 9694 99 9728 133
rect 9762 99 9796 133
rect 9830 99 9864 133
rect 9898 99 9932 133
rect 9966 99 10000 133
rect 10034 99 10068 133
rect 10102 99 10136 133
rect 10170 99 10204 133
rect 10238 99 10272 133
rect 10306 99 10340 133
rect 10374 99 10408 133
rect 10442 99 10476 133
rect 10510 99 10544 133
rect 10578 99 10612 133
rect 10646 99 10680 133
rect 10714 99 10748 133
rect 10782 99 10816 133
rect 10850 99 10884 133
rect 10918 99 10952 133
rect 10986 99 11020 133
rect 11054 99 11088 133
rect 11122 99 11156 133
rect 11190 99 11224 133
rect 11258 99 11292 133
rect 11326 99 11360 133
rect 11394 99 11428 133
rect 11462 99 11496 133
rect 11530 99 11564 133
rect 11598 99 11632 133
rect 11666 99 11700 133
rect 11734 99 11768 133
rect 11802 99 11836 133
rect 11870 99 11904 133
rect 11938 99 11972 133
rect 12006 99 12040 133
rect 12074 99 12098 133
rect 1719 61 1889 95
rect 1048 -30 1110 34
rect 1313 -15 1889 61
rect 1313 -49 1783 -15
rect 1817 -49 1855 -15
rect 3030 -7 3275 17
rect 3064 -41 3136 -7
rect 3170 -41 3241 -7
rect 3030 -65 3275 -41
rect 4583 -25 4689 61
rect 4617 -59 4655 -25
rect 1340 -124 1573 -120
rect 1607 -124 1646 -119
rect 1680 -124 1719 -119
rect 1753 -124 1792 -119
rect 1826 -124 1865 -119
rect 1899 -124 1938 -119
rect 1972 -124 2011 -119
rect 2045 -124 2084 -119
rect 2118 -124 2157 -119
rect 2191 -124 2230 -119
rect 2264 -124 2303 -119
rect 2337 -124 2376 -119
rect 2410 -124 2449 -119
rect 2483 -124 2522 -119
rect 2556 -124 2595 -119
rect 2629 -124 2668 -119
rect 2702 -124 2741 -119
rect 1340 -158 1374 -124
rect 1408 -158 1445 -124
rect 1479 -158 1516 -124
rect 1550 -153 1573 -124
rect 1621 -153 1646 -124
rect 1691 -153 1719 -124
rect 1761 -153 1792 -124
rect 1831 -153 1865 -124
rect 1550 -158 1587 -153
rect 1621 -158 1657 -153
rect 1691 -158 1727 -153
rect 1761 -158 1797 -153
rect 1831 -158 1867 -153
rect 1901 -158 1937 -124
rect 1972 -153 2007 -124
rect 2045 -153 2077 -124
rect 2118 -153 2147 -124
rect 2191 -153 2217 -124
rect 2264 -153 2287 -124
rect 2337 -153 2357 -124
rect 2410 -153 2427 -124
rect 2483 -153 2497 -124
rect 2556 -153 2567 -124
rect 2629 -153 2637 -124
rect 2702 -153 2707 -124
rect 1971 -158 2007 -153
rect 2041 -158 2077 -153
rect 2111 -158 2147 -153
rect 2181 -158 2217 -153
rect 2251 -158 2287 -153
rect 2321 -158 2357 -153
rect 2391 -158 2427 -153
rect 2461 -158 2497 -153
rect 2531 -158 2567 -153
rect 2601 -158 2637 -153
rect 2671 -158 2707 -153
rect 2775 -124 2814 -119
rect 2848 -124 2887 -119
rect 2921 -124 2960 -119
rect 2994 -124 3033 -119
rect 3067 -124 3106 -119
rect 3140 -124 3179 -119
rect 3213 -124 3252 -119
rect 3286 -124 3325 -119
rect 3359 -124 3398 -119
rect 3432 -124 3471 -119
rect 3505 -124 3544 -119
rect 3578 -124 3617 -119
rect 2775 -153 2777 -124
rect 2741 -158 2777 -153
rect 2811 -153 2814 -124
rect 2881 -153 2887 -124
rect 2951 -153 2960 -124
rect 3021 -153 3033 -124
rect 3091 -153 3106 -124
rect 3161 -153 3179 -124
rect 3231 -153 3252 -124
rect 3301 -153 3325 -124
rect 3371 -153 3398 -124
rect 3441 -153 3471 -124
rect 3511 -153 3544 -124
rect 2811 -158 2847 -153
rect 2881 -158 2917 -153
rect 2951 -158 2987 -153
rect 3021 -158 3057 -153
rect 3091 -158 3127 -153
rect 3161 -158 3197 -153
rect 3231 -158 3267 -153
rect 3301 -158 3337 -153
rect 3371 -158 3407 -153
rect 3441 -158 3477 -153
rect 3511 -158 3547 -153
rect 3581 -158 3617 -124
rect 3651 -153 3690 -119
rect 3724 -153 3763 -119
rect 3797 -153 3836 -119
rect 3870 -153 3909 -119
rect 3943 -153 3982 -119
rect 4016 -153 4055 -119
rect 4089 -153 4128 -119
rect 4162 -153 4201 -119
rect 4235 -153 4274 -119
rect 4308 -153 4347 -119
rect 4381 -153 4420 -119
rect 4454 -153 4493 -119
rect 4527 -153 4565 -119
rect 4599 -153 4637 -119
rect 4671 -153 4709 -119
rect 3651 -158 4743 -153
rect 1340 -194 4743 -158
rect 1340 -228 1374 -194
rect 1408 -228 1445 -194
rect 1479 -228 1516 -194
rect 1550 -201 1587 -194
rect 1621 -201 1657 -194
rect 1691 -201 1727 -194
rect 1761 -201 1797 -194
rect 1831 -201 1867 -194
rect 1550 -228 1573 -201
rect 1621 -228 1646 -201
rect 1691 -228 1719 -201
rect 1761 -228 1792 -201
rect 1831 -228 1865 -201
rect 1901 -228 1937 -194
rect 1971 -201 2007 -194
rect 2041 -201 2077 -194
rect 2111 -201 2147 -194
rect 2181 -201 2217 -194
rect 2251 -201 2287 -194
rect 2321 -201 2357 -194
rect 2391 -201 2427 -194
rect 2461 -201 2497 -194
rect 2531 -201 2567 -194
rect 2601 -201 2637 -194
rect 2671 -201 2707 -194
rect 1972 -228 2007 -201
rect 2045 -228 2077 -201
rect 2118 -228 2147 -201
rect 2191 -228 2217 -201
rect 2264 -228 2287 -201
rect 2337 -228 2357 -201
rect 2410 -228 2427 -201
rect 2483 -228 2497 -201
rect 2556 -228 2567 -201
rect 2629 -228 2637 -201
rect 2702 -228 2707 -201
rect 2741 -201 2777 -194
rect 1340 -235 1573 -228
rect 1607 -235 1646 -228
rect 1680 -235 1719 -228
rect 1753 -235 1792 -228
rect 1826 -235 1865 -228
rect 1899 -235 1938 -228
rect 1972 -235 2011 -228
rect 2045 -235 2084 -228
rect 2118 -235 2157 -228
rect 2191 -235 2230 -228
rect 2264 -235 2303 -228
rect 2337 -235 2376 -228
rect 2410 -235 2449 -228
rect 2483 -235 2522 -228
rect 2556 -235 2595 -228
rect 2629 -235 2668 -228
rect 2702 -235 2741 -228
rect 2775 -228 2777 -201
rect 2811 -201 2847 -194
rect 2881 -201 2917 -194
rect 2951 -201 2987 -194
rect 3021 -201 3057 -194
rect 3091 -201 3127 -194
rect 3161 -201 3197 -194
rect 3231 -201 3267 -194
rect 3301 -201 3337 -194
rect 3371 -201 3407 -194
rect 3441 -201 3477 -194
rect 3511 -201 3547 -194
rect 2811 -228 2814 -201
rect 2881 -228 2887 -201
rect 2951 -228 2960 -201
rect 3021 -228 3033 -201
rect 3091 -228 3106 -201
rect 3161 -228 3179 -201
rect 3231 -228 3252 -201
rect 3301 -228 3325 -201
rect 3371 -228 3398 -201
rect 3441 -228 3471 -201
rect 3511 -228 3544 -201
rect 3581 -228 3617 -194
rect 3651 -201 4743 -194
rect 2775 -235 2814 -228
rect 2848 -235 2887 -228
rect 2921 -235 2960 -228
rect 2994 -235 3033 -228
rect 3067 -235 3106 -228
rect 3140 -235 3179 -228
rect 3213 -235 3252 -228
rect 3286 -235 3325 -228
rect 3359 -235 3398 -228
rect 3432 -235 3471 -228
rect 3505 -235 3544 -228
rect 3578 -235 3617 -228
rect 3651 -235 3690 -201
rect 3724 -235 3763 -201
rect 3797 -235 3836 -201
rect 3870 -235 3909 -201
rect 3943 -235 3982 -201
rect 4016 -235 4055 -201
rect 4089 -235 4128 -201
rect 4162 -235 4201 -201
rect 4235 -235 4274 -201
rect 4308 -235 4347 -201
rect 4381 -235 4420 -201
rect 4454 -235 4493 -201
rect 4527 -235 4565 -201
rect 4599 -235 4637 -201
rect 4671 -235 4709 -201
rect 1340 -264 3685 -235
rect 1340 -298 1374 -264
rect 1408 -298 1445 -264
rect 1479 -298 1516 -264
rect 1550 -298 1587 -264
rect 1621 -298 1657 -264
rect 1691 -298 1727 -264
rect 1761 -298 1797 -264
rect 1831 -298 1867 -264
rect 1901 -298 1937 -264
rect 1971 -298 2007 -264
rect 2041 -298 2077 -264
rect 2111 -298 2147 -264
rect 2181 -298 2217 -264
rect 2251 -298 2287 -264
rect 2321 -298 2357 -264
rect 2391 -298 2427 -264
rect 2461 -298 2497 -264
rect 2531 -298 2567 -264
rect 2601 -298 2637 -264
rect 2671 -298 2707 -264
rect 2741 -298 2777 -264
rect 2811 -298 2847 -264
rect 2881 -298 2917 -264
rect 2951 -298 2987 -264
rect 3021 -298 3057 -264
rect 3091 -298 3127 -264
rect 3161 -298 3197 -264
rect 3231 -298 3267 -264
rect 3301 -298 3337 -264
rect 3371 -298 3407 -264
rect 3441 -298 3477 -264
rect 3511 -298 3547 -264
rect 3581 -298 3617 -264
rect 3651 -298 3685 -264
rect 1340 -308 3685 -298
rect -227 -313 3685 -308
rect -227 -347 -193 -313
rect -159 -347 -123 -313
rect -89 -347 -53 -313
rect -19 -347 17 -313
rect 51 -347 87 -313
rect 121 -347 157 -313
rect 191 -347 227 -313
rect 261 -347 297 -313
rect 331 -347 367 -313
rect 401 -347 437 -313
rect 471 -347 507 -313
rect 541 -347 577 -313
rect 611 -347 647 -313
rect 681 -347 717 -313
rect 751 -347 787 -313
rect 821 -347 857 -313
rect 891 -347 927 -313
rect 961 -347 996 -313
rect 1030 -347 1065 -313
rect 1099 -347 1134 -313
rect 1168 -347 1203 -313
rect 1237 -347 1272 -313
rect 1306 -334 3685 -313
rect 1306 -347 1374 -334
rect -227 -368 1374 -347
rect 1408 -368 1445 -334
rect 1479 -368 1516 -334
rect 1550 -368 1587 -334
rect 1621 -368 1657 -334
rect 1691 -368 1727 -334
rect 1761 -368 1797 -334
rect 1831 -368 1867 -334
rect 1901 -368 1937 -334
rect 1971 -368 2007 -334
rect 2041 -368 2077 -334
rect 2111 -368 2147 -334
rect 2181 -368 2217 -334
rect 2251 -368 2287 -334
rect 2321 -368 2357 -334
rect 2391 -368 2427 -334
rect 2461 -368 2497 -334
rect 2531 -368 2567 -334
rect 2601 -368 2637 -334
rect 2671 -368 2707 -334
rect 2741 -368 2777 -334
rect 2811 -368 2847 -334
rect 2881 -368 2917 -334
rect 2951 -368 2987 -334
rect 3021 -368 3057 -334
rect 3091 -368 3127 -334
rect 3161 -368 3197 -334
rect 3231 -368 3267 -334
rect 3301 -368 3337 -334
rect 3371 -368 3407 -334
rect 3441 -368 3477 -334
rect 3511 -368 3547 -334
rect 3581 -368 3617 -334
rect 3651 -368 3685 -334
rect -227 -385 3685 -368
rect -227 -419 -193 -385
rect -159 -419 -123 -385
rect -89 -419 -53 -385
rect -19 -419 17 -385
rect 51 -419 87 -385
rect 121 -419 157 -385
rect 191 -419 227 -385
rect 261 -419 297 -385
rect 331 -419 367 -385
rect 401 -419 437 -385
rect 471 -419 507 -385
rect 541 -419 577 -385
rect 611 -419 647 -385
rect 681 -419 717 -385
rect 751 -419 787 -385
rect 821 -419 857 -385
rect 891 -419 927 -385
rect 961 -419 996 -385
rect 1030 -419 1065 -385
rect 1099 -419 1134 -385
rect 1168 -419 1203 -385
rect 1237 -419 1272 -385
rect 1306 -404 3685 -385
rect 1306 -419 1374 -404
rect -227 -438 1374 -419
rect 1408 -438 1445 -404
rect 1479 -438 1516 -404
rect 1550 -438 1587 -404
rect 1621 -438 1657 -404
rect 1691 -438 1727 -404
rect 1761 -438 1797 -404
rect 1831 -438 1867 -404
rect 1901 -438 1937 -404
rect 1971 -438 2007 -404
rect 2041 -438 2077 -404
rect 2111 -438 2147 -404
rect 2181 -438 2217 -404
rect 2251 -438 2287 -404
rect 2321 -438 2357 -404
rect 2391 -438 2427 -404
rect 2461 -438 2497 -404
rect 2531 -438 2567 -404
rect 2601 -438 2637 -404
rect 2671 -438 2707 -404
rect 2741 -438 2777 -404
rect 2811 -438 2847 -404
rect 2881 -438 2917 -404
rect 2951 -438 2987 -404
rect 3021 -438 3057 -404
rect 3091 -438 3127 -404
rect 3161 -438 3197 -404
rect 3231 -438 3267 -404
rect 3301 -438 3337 -404
rect 3371 -438 3407 -404
rect 3441 -438 3477 -404
rect 3511 -438 3547 -404
rect 3581 -438 3617 -404
rect 3651 -438 3685 -404
rect -227 -457 3685 -438
rect -227 -491 -193 -457
rect -159 -491 -123 -457
rect -89 -491 -53 -457
rect -19 -491 17 -457
rect 51 -491 87 -457
rect 121 -491 157 -457
rect 191 -491 227 -457
rect 261 -491 297 -457
rect 331 -491 367 -457
rect 401 -491 437 -457
rect 471 -491 507 -457
rect 541 -491 577 -457
rect 611 -491 647 -457
rect 681 -491 717 -457
rect 751 -491 787 -457
rect 821 -491 857 -457
rect 891 -491 927 -457
rect 961 -491 996 -457
rect 1030 -491 1065 -457
rect 1099 -491 1134 -457
rect 1168 -491 1203 -457
rect 1237 -491 1272 -457
rect 1306 -474 3685 -457
rect 1306 -491 1374 -474
rect -227 -508 1374 -491
rect 1408 -508 1445 -474
rect 1479 -508 1516 -474
rect 1550 -508 1587 -474
rect 1621 -508 1657 -474
rect 1691 -508 1727 -474
rect 1761 -508 1797 -474
rect 1831 -508 1867 -474
rect 1901 -508 1937 -474
rect 1971 -508 2007 -474
rect 2041 -508 2077 -474
rect 2111 -508 2147 -474
rect 2181 -508 2217 -474
rect 2251 -508 2287 -474
rect 2321 -508 2357 -474
rect 2391 -508 2427 -474
rect 2461 -508 2497 -474
rect 2531 -508 2567 -474
rect 2601 -508 2637 -474
rect 2671 -508 2707 -474
rect 2741 -508 2777 -474
rect 2811 -508 2847 -474
rect 2881 -508 2917 -474
rect 2951 -508 2987 -474
rect 3021 -508 3057 -474
rect 3091 -508 3127 -474
rect 3161 -508 3197 -474
rect 3231 -508 3267 -474
rect 3301 -508 3337 -474
rect 3371 -508 3407 -474
rect 3441 -508 3477 -474
rect 3511 -508 3547 -474
rect 3581 -508 3617 -474
rect 3651 -508 3685 -474
rect -227 -529 3685 -508
rect -227 -563 -193 -529
rect -159 -563 -123 -529
rect -89 -563 -53 -529
rect -19 -563 17 -529
rect 51 -563 87 -529
rect 121 -563 157 -529
rect 191 -563 227 -529
rect 261 -563 297 -529
rect 331 -563 367 -529
rect 401 -563 437 -529
rect 471 -563 507 -529
rect 541 -563 577 -529
rect 611 -563 647 -529
rect 681 -563 717 -529
rect 751 -563 787 -529
rect 821 -563 857 -529
rect 891 -563 927 -529
rect 961 -563 996 -529
rect 1030 -563 1065 -529
rect 1099 -563 1134 -529
rect 1168 -563 1203 -529
rect 1237 -563 1272 -529
rect 1306 -544 3685 -529
rect 1306 -563 1374 -544
rect -227 -578 1374 -563
rect 1408 -578 1445 -544
rect 1479 -578 1516 -544
rect 1550 -578 1587 -544
rect 1621 -578 1657 -544
rect 1691 -578 1727 -544
rect 1761 -578 1797 -544
rect 1831 -578 1867 -544
rect 1901 -578 1937 -544
rect 1971 -578 2007 -544
rect 2041 -578 2077 -544
rect 2111 -578 2147 -544
rect 2181 -578 2217 -544
rect 2251 -578 2287 -544
rect 2321 -578 2357 -544
rect 2391 -578 2427 -544
rect 2461 -578 2497 -544
rect 2531 -578 2567 -544
rect 2601 -578 2637 -544
rect 2671 -578 2707 -544
rect 2741 -578 2777 -544
rect 2811 -578 2847 -544
rect 2881 -578 2917 -544
rect 2951 -578 2987 -544
rect 3021 -578 3057 -544
rect 3091 -578 3127 -544
rect 3161 -578 3197 -544
rect 3231 -578 3267 -544
rect 3301 -578 3337 -544
rect 3371 -578 3407 -544
rect 3441 -578 3477 -544
rect 3511 -578 3547 -544
rect 3581 -578 3617 -544
rect 3651 -578 3685 -544
rect -227 -601 3685 -578
rect -227 -635 -193 -601
rect -159 -635 -123 -601
rect -89 -635 -53 -601
rect -19 -635 17 -601
rect 51 -635 87 -601
rect 121 -635 157 -601
rect 191 -635 227 -601
rect 261 -635 297 -601
rect 331 -635 367 -601
rect 401 -635 437 -601
rect 471 -635 507 -601
rect 541 -635 577 -601
rect 611 -635 647 -601
rect 681 -635 717 -601
rect 751 -635 787 -601
rect 821 -635 857 -601
rect 891 -635 927 -601
rect 961 -635 996 -601
rect 1030 -635 1065 -601
rect 1099 -635 1134 -601
rect 1168 -635 1203 -601
rect 1237 -635 1272 -601
rect 1306 -614 3685 -601
rect 1306 -635 1374 -614
rect -227 -648 1374 -635
rect 1408 -648 1445 -614
rect 1479 -648 1516 -614
rect 1550 -648 1587 -614
rect 1621 -648 1657 -614
rect 1691 -648 1727 -614
rect 1761 -648 1797 -614
rect 1831 -648 1867 -614
rect 1901 -648 1937 -614
rect 1971 -648 2007 -614
rect 2041 -648 2077 -614
rect 2111 -648 2147 -614
rect 2181 -648 2217 -614
rect 2251 -648 2287 -614
rect 2321 -648 2357 -614
rect 2391 -648 2427 -614
rect 2461 -648 2497 -614
rect 2531 -648 2567 -614
rect 2601 -648 2637 -614
rect 2671 -648 2707 -614
rect 2741 -648 2777 -614
rect 2811 -648 2847 -614
rect 2881 -648 2917 -614
rect 2951 -648 2987 -614
rect 3021 -648 3057 -614
rect 3091 -648 3127 -614
rect 3161 -648 3197 -614
rect 3231 -648 3267 -614
rect 3301 -648 3337 -614
rect 3371 -648 3407 -614
rect 3441 -648 3477 -614
rect 3511 -648 3547 -614
rect 3581 -648 3617 -614
rect 3651 -648 3685 -614
rect -227 -673 3685 -648
rect -227 -707 -193 -673
rect -159 -707 -123 -673
rect -89 -707 -53 -673
rect -19 -707 17 -673
rect 51 -707 87 -673
rect 121 -707 157 -673
rect 191 -707 227 -673
rect 261 -707 297 -673
rect 331 -707 367 -673
rect 401 -707 437 -673
rect 471 -707 507 -673
rect 541 -707 577 -673
rect 611 -707 647 -673
rect 681 -707 717 -673
rect 751 -707 787 -673
rect 821 -707 857 -673
rect 891 -707 927 -673
rect 961 -707 996 -673
rect 1030 -707 1065 -673
rect 1099 -707 1134 -673
rect 1168 -707 1203 -673
rect 1237 -707 1272 -673
rect 1306 -684 3685 -673
rect 1306 -707 1374 -684
rect -227 -718 1374 -707
rect 1408 -718 1445 -684
rect 1479 -718 1516 -684
rect 1550 -718 1587 -684
rect 1621 -718 1657 -684
rect 1691 -718 1727 -684
rect 1761 -718 1797 -684
rect 1831 -718 1867 -684
rect 1901 -718 1937 -684
rect 1971 -718 2007 -684
rect 2041 -718 2077 -684
rect 2111 -718 2147 -684
rect 2181 -718 2217 -684
rect 2251 -718 2287 -684
rect 2321 -718 2357 -684
rect 2391 -718 2427 -684
rect 2461 -718 2497 -684
rect 2531 -718 2567 -684
rect 2601 -718 2637 -684
rect 2671 -718 2707 -684
rect 2741 -718 2777 -684
rect 2811 -718 2847 -684
rect 2881 -718 2917 -684
rect 2951 -718 2987 -684
rect 3021 -718 3057 -684
rect 3091 -718 3127 -684
rect 3161 -718 3197 -684
rect 3231 -718 3267 -684
rect 3301 -718 3337 -684
rect 3371 -718 3407 -684
rect 3441 -718 3477 -684
rect 3511 -718 3547 -684
rect 3581 -718 3617 -684
rect 3651 -718 3685 -684
rect -227 -745 3685 -718
rect -227 -779 -193 -745
rect -159 -779 -123 -745
rect -89 -779 -53 -745
rect -19 -779 17 -745
rect 51 -779 87 -745
rect 121 -779 157 -745
rect 191 -779 227 -745
rect 261 -779 297 -745
rect 331 -779 367 -745
rect 401 -779 437 -745
rect 471 -779 507 -745
rect 541 -779 577 -745
rect 611 -779 647 -745
rect 681 -779 717 -745
rect 751 -779 787 -745
rect 821 -779 857 -745
rect 891 -779 927 -745
rect 961 -779 996 -745
rect 1030 -779 1065 -745
rect 1099 -779 1134 -745
rect 1168 -779 1203 -745
rect 1237 -779 1272 -745
rect 1306 -754 3685 -745
rect 1306 -779 1374 -754
rect -227 -788 1374 -779
rect 1408 -788 1445 -754
rect 1479 -788 1516 -754
rect 1550 -788 1587 -754
rect 1621 -788 1657 -754
rect 1691 -788 1727 -754
rect 1761 -788 1797 -754
rect 1831 -788 1867 -754
rect 1901 -788 1937 -754
rect 1971 -788 2007 -754
rect 2041 -788 2077 -754
rect 2111 -788 2147 -754
rect 2181 -788 2217 -754
rect 2251 -788 2287 -754
rect 2321 -788 2357 -754
rect 2391 -788 2427 -754
rect 2461 -788 2497 -754
rect 2531 -788 2567 -754
rect 2601 -788 2637 -754
rect 2671 -788 2707 -754
rect 2741 -788 2777 -754
rect 2811 -788 2847 -754
rect 2881 -788 2917 -754
rect 2951 -788 2987 -754
rect 3021 -788 3057 -754
rect 3091 -788 3127 -754
rect 3161 -788 3197 -754
rect 3231 -788 3267 -754
rect 3301 -788 3337 -754
rect 3371 -788 3407 -754
rect 3441 -788 3477 -754
rect 3511 -788 3547 -754
rect 3581 -788 3617 -754
rect 3651 -788 3685 -754
rect -227 -817 3685 -788
rect -227 -851 -193 -817
rect -159 -851 -123 -817
rect -89 -851 -53 -817
rect -19 -851 17 -817
rect 51 -851 87 -817
rect 121 -851 157 -817
rect 191 -851 227 -817
rect 261 -851 297 -817
rect 331 -851 367 -817
rect 401 -851 437 -817
rect 471 -851 507 -817
rect 541 -851 577 -817
rect 611 -851 647 -817
rect 681 -851 717 -817
rect 751 -851 787 -817
rect 821 -851 857 -817
rect 891 -851 927 -817
rect 961 -851 996 -817
rect 1030 -851 1065 -817
rect 1099 -851 1134 -817
rect 1168 -851 1203 -817
rect 1237 -851 1272 -817
rect 1306 -824 3685 -817
rect 1306 -851 1374 -824
rect -227 -858 1374 -851
rect 1408 -858 1445 -824
rect 1479 -858 1516 -824
rect 1550 -858 1587 -824
rect 1621 -858 1657 -824
rect 1691 -858 1727 -824
rect 1761 -858 1797 -824
rect 1831 -858 1867 -824
rect 1901 -858 1937 -824
rect 1971 -858 2007 -824
rect 2041 -858 2077 -824
rect 2111 -858 2147 -824
rect 2181 -858 2217 -824
rect 2251 -858 2287 -824
rect 2321 -858 2357 -824
rect 2391 -858 2427 -824
rect 2461 -858 2497 -824
rect 2531 -858 2567 -824
rect 2601 -858 2637 -824
rect 2671 -858 2707 -824
rect 2741 -858 2777 -824
rect 2811 -858 2847 -824
rect 2881 -858 2917 -824
rect 2951 -858 2987 -824
rect 3021 -858 3057 -824
rect 3091 -858 3127 -824
rect 3161 -858 3197 -824
rect 3231 -858 3267 -824
rect 3301 -858 3337 -824
rect 3371 -858 3407 -824
rect 3441 -858 3477 -824
rect 3511 -858 3547 -824
rect 3581 -858 3617 -824
rect 3651 -858 3685 -824
rect -227 -889 3685 -858
rect -227 -923 -193 -889
rect -159 -923 -123 -889
rect -89 -923 -53 -889
rect -19 -923 17 -889
rect 51 -923 87 -889
rect 121 -923 157 -889
rect 191 -923 227 -889
rect 261 -923 297 -889
rect 331 -923 367 -889
rect 401 -923 437 -889
rect 471 -923 507 -889
rect 541 -923 577 -889
rect 611 -923 647 -889
rect 681 -923 717 -889
rect 751 -923 787 -889
rect 821 -923 857 -889
rect 891 -923 927 -889
rect 961 -923 996 -889
rect 1030 -923 1065 -889
rect 1099 -923 1134 -889
rect 1168 -923 1203 -889
rect 1237 -923 1272 -889
rect 1306 -894 3685 -889
rect 1306 -923 1374 -894
rect -227 -928 1374 -923
rect 1408 -928 1445 -894
rect 1479 -912 1516 -894
rect 1479 -928 1480 -912
rect -227 -946 1480 -928
rect 1514 -928 1516 -912
rect 1550 -912 1587 -894
rect 1621 -912 1657 -894
rect 1691 -912 1727 -894
rect 1761 -912 1797 -894
rect 1831 -912 1867 -894
rect 1901 -912 1937 -894
rect 1550 -928 1556 -912
rect 1621 -928 1632 -912
rect 1691 -928 1707 -912
rect 1761 -928 1782 -912
rect 1831 -928 1857 -912
rect 1901 -928 1932 -912
rect 1971 -928 2007 -894
rect 2041 -928 2077 -894
rect 2111 -912 2147 -894
rect 2181 -912 2217 -894
rect 2251 -912 2287 -894
rect 2321 -912 2357 -894
rect 2391 -912 2427 -894
rect 2461 -912 2497 -894
rect 2116 -928 2147 -912
rect 2191 -928 2217 -912
rect 2266 -928 2287 -912
rect 2341 -928 2357 -912
rect 2416 -928 2427 -912
rect 2491 -928 2497 -912
rect 2531 -912 2567 -894
rect 2531 -928 2532 -912
rect 1514 -946 1556 -928
rect 1590 -946 1632 -928
rect 1666 -946 1707 -928
rect 1741 -946 1782 -928
rect 1816 -946 1857 -928
rect 1891 -946 1932 -928
rect 1966 -946 2007 -928
rect 2041 -946 2082 -928
rect 2116 -946 2157 -928
rect 2191 -946 2232 -928
rect 2266 -946 2307 -928
rect 2341 -946 2382 -928
rect 2416 -946 2457 -928
rect 2491 -946 2532 -928
rect 2566 -928 2567 -912
rect 2601 -912 2637 -894
rect 2671 -912 2707 -894
rect 2741 -912 2777 -894
rect 2811 -912 2847 -894
rect 2881 -912 2917 -894
rect 2951 -912 2987 -894
rect 2601 -928 2607 -912
rect 2671 -928 2682 -912
rect 2741 -928 2757 -912
rect 2811 -928 2832 -912
rect 2881 -928 2907 -912
rect 2951 -928 2982 -912
rect 3021 -928 3057 -894
rect 3091 -928 3127 -894
rect 3161 -912 3197 -894
rect 3231 -912 3267 -894
rect 3166 -928 3197 -912
rect 3241 -928 3267 -912
rect 3301 -928 3337 -894
rect 3371 -928 3407 -894
rect 3441 -928 3477 -894
rect 3511 -928 3547 -894
rect 3581 -928 3617 -894
rect 3651 -928 3685 -894
rect 2566 -946 2607 -928
rect 2641 -946 2682 -928
rect 2716 -946 2757 -928
rect 2791 -946 2832 -928
rect 2866 -946 2907 -928
rect 2941 -946 2982 -928
rect 3016 -946 3057 -928
rect 3091 -946 3132 -928
rect 3166 -946 3207 -928
rect 3241 -946 3685 -928
rect -227 -961 3685 -946
rect -227 -995 -193 -961
rect -159 -995 -123 -961
rect -89 -995 -53 -961
rect -19 -995 17 -961
rect 51 -995 87 -961
rect 121 -995 157 -961
rect 191 -995 227 -961
rect 261 -995 297 -961
rect 331 -995 367 -961
rect 401 -995 437 -961
rect 471 -995 507 -961
rect 541 -995 577 -961
rect 611 -995 647 -961
rect 681 -995 717 -961
rect 751 -995 787 -961
rect 821 -995 857 -961
rect 891 -995 927 -961
rect 961 -995 996 -961
rect 1030 -995 1065 -961
rect 1099 -995 1134 -961
rect 1168 -995 1203 -961
rect 1237 -995 1272 -961
rect 1306 -964 3685 -961
rect 1306 -995 1374 -964
rect -227 -998 1374 -995
rect 1408 -998 1445 -964
rect 1479 -998 1516 -964
rect 1550 -998 1587 -964
rect 1621 -998 1657 -964
rect 1691 -998 1727 -964
rect 1761 -998 1797 -964
rect 1831 -998 1867 -964
rect 1901 -998 1937 -964
rect 1971 -998 2007 -964
rect 2041 -998 2077 -964
rect 2111 -998 2147 -964
rect 2181 -998 2217 -964
rect 2251 -998 2287 -964
rect 2321 -998 2357 -964
rect 2391 -998 2427 -964
rect 2461 -998 2497 -964
rect 2531 -998 2567 -964
rect 2601 -998 2637 -964
rect 2671 -998 2707 -964
rect 2741 -998 2777 -964
rect 2811 -998 2847 -964
rect 2881 -998 2917 -964
rect 2951 -998 2987 -964
rect 3021 -998 3057 -964
rect 3091 -998 3127 -964
rect 3161 -998 3197 -964
rect 3231 -998 3267 -964
rect 3301 -998 3337 -964
rect 3371 -998 3407 -964
rect 3441 -998 3477 -964
rect 3511 -998 3547 -964
rect 3581 -998 3617 -964
rect 3651 -998 3685 -964
rect -227 -1033 3685 -998
rect -227 -1067 -193 -1033
rect -159 -1067 -123 -1033
rect -89 -1067 -53 -1033
rect -19 -1067 17 -1033
rect 51 -1067 87 -1033
rect 121 -1067 157 -1033
rect 191 -1067 227 -1033
rect 261 -1067 297 -1033
rect 331 -1067 367 -1033
rect 401 -1067 437 -1033
rect 471 -1067 507 -1033
rect 541 -1067 577 -1033
rect 611 -1067 647 -1033
rect 681 -1067 717 -1033
rect 751 -1067 787 -1033
rect 821 -1067 857 -1033
rect 891 -1067 927 -1033
rect 961 -1067 996 -1033
rect 1030 -1067 1065 -1033
rect 1099 -1067 1134 -1033
rect 1168 -1067 1203 -1033
rect 1237 -1067 1272 -1033
rect 1306 -1034 3685 -1033
rect 1306 -1067 1374 -1034
rect -227 -1068 1374 -1067
rect 1408 -1068 1445 -1034
rect 1479 -1068 1516 -1034
rect 1550 -1068 1587 -1034
rect 1621 -1068 1657 -1034
rect 1691 -1068 1727 -1034
rect 1761 -1068 1797 -1034
rect 1831 -1068 1867 -1034
rect 1901 -1068 1937 -1034
rect 1971 -1068 2007 -1034
rect 2041 -1068 2077 -1034
rect 2111 -1068 2147 -1034
rect 2181 -1068 2217 -1034
rect 2251 -1068 2287 -1034
rect 2321 -1068 2357 -1034
rect 2391 -1068 2427 -1034
rect 2461 -1068 2497 -1034
rect 2531 -1068 2567 -1034
rect 2601 -1068 2637 -1034
rect 2671 -1068 2707 -1034
rect 2741 -1068 2777 -1034
rect 2811 -1068 2847 -1034
rect 2881 -1068 2917 -1034
rect 2951 -1068 2987 -1034
rect 3021 -1068 3057 -1034
rect 3091 -1068 3127 -1034
rect 3161 -1068 3197 -1034
rect 3231 -1068 3267 -1034
rect 3301 -1068 3337 -1034
rect 3371 -1068 3407 -1034
rect 3441 -1068 3477 -1034
rect 3511 -1068 3547 -1034
rect 3581 -1068 3617 -1034
rect 3651 -1068 3685 -1034
rect -227 -1072 3685 -1068
<< viali >>
rect 2582 1967 2596 1999
rect 2596 1967 2616 1999
rect 2655 1967 2669 1999
rect 2669 1967 2689 1999
rect 2728 1967 2741 1999
rect 2741 1967 2762 1999
rect 2801 1967 2813 1999
rect 2813 1967 2835 1999
rect 2874 1967 2885 1999
rect 2885 1967 2908 1999
rect 2947 1967 2957 1999
rect 2957 1967 2981 1999
rect 3020 1967 3029 1999
rect 3029 1967 3054 1999
rect 3092 1967 3101 1999
rect 3101 1967 3126 1999
rect 3164 1967 3173 1999
rect 3173 1967 3198 1999
rect 3236 1967 3245 1999
rect 3245 1967 3270 1999
rect 3308 1967 3317 1999
rect 3317 1967 3342 1999
rect 3380 1967 3389 1999
rect 3389 1967 3414 1999
rect 3452 1967 3461 1999
rect 3461 1967 3486 1999
rect 3524 1967 3533 1999
rect 3533 1967 3558 1999
rect 3596 1967 3605 1999
rect 3605 1967 3630 1999
rect 3668 1967 3677 1999
rect 3677 1967 3702 1999
rect 2582 1965 2616 1967
rect 2655 1965 2689 1967
rect 2728 1965 2762 1967
rect 2801 1965 2835 1967
rect 2874 1965 2908 1967
rect 2947 1965 2981 1967
rect 3020 1965 3054 1967
rect 3092 1965 3126 1967
rect 3164 1965 3198 1967
rect 3236 1965 3270 1967
rect 3308 1965 3342 1967
rect 3380 1965 3414 1967
rect 3452 1965 3486 1967
rect 3524 1965 3558 1967
rect 3596 1965 3630 1967
rect 3668 1965 3702 1967
rect 2582 1899 2613 1915
rect 2613 1899 2616 1915
rect 2655 1899 2682 1915
rect 2682 1899 2689 1915
rect 2728 1899 2751 1915
rect 2751 1899 2762 1915
rect 2801 1899 2820 1915
rect 2820 1899 2835 1915
rect 2874 1899 2889 1915
rect 2889 1899 2908 1915
rect 2947 1899 2958 1915
rect 2958 1899 2981 1915
rect 3020 1899 3027 1915
rect 3027 1899 3054 1915
rect 3092 1899 3096 1915
rect 3096 1899 3126 1915
rect 3164 1899 3165 1915
rect 3165 1899 3198 1915
rect 3236 1899 3269 1915
rect 3269 1899 3270 1915
rect 3308 1899 3338 1915
rect 3338 1899 3342 1915
rect 3380 1899 3407 1915
rect 3407 1899 3414 1915
rect 3452 1899 3476 1915
rect 3476 1899 3486 1915
rect 3524 1899 3545 1915
rect 3545 1899 3558 1915
rect 3596 1899 3613 1915
rect 3613 1899 3630 1915
rect 3668 1899 3681 1915
rect 3681 1899 3702 1915
rect 2582 1881 2616 1899
rect 2655 1881 2689 1899
rect 2728 1881 2762 1899
rect 2801 1881 2835 1899
rect 2874 1881 2908 1899
rect 2947 1881 2981 1899
rect 3020 1881 3054 1899
rect 3092 1881 3126 1899
rect 3164 1881 3198 1899
rect 3236 1881 3270 1899
rect 3308 1881 3342 1899
rect 3380 1881 3414 1899
rect 3452 1881 3486 1899
rect 3524 1881 3558 1899
rect 3596 1881 3630 1899
rect 3668 1881 3702 1899
rect 488 1549 522 1583
rect 560 1549 594 1583
rect 5797 1167 5831 1201
rect 5869 1167 5903 1201
rect 11785 1107 12323 1213
rect 868 1018 902 1052
rect 868 946 902 980
rect 5218 590 5252 624
rect 5218 518 5252 552
rect 5394 1006 5428 1040
rect 7050 1040 7084 1074
rect 7050 968 7084 1002
rect 5394 934 5428 968
rect 1783 -49 1817 -15
rect 1855 -49 1889 -15
rect 3030 -41 3064 -7
rect 3136 -41 3170 -7
rect 3241 -41 3275 -7
rect 4583 -59 4617 -25
rect 4655 -59 4689 -25
rect 1573 -124 1607 -119
rect 1646 -124 1680 -119
rect 1719 -124 1753 -119
rect 1792 -124 1826 -119
rect 1865 -124 1899 -119
rect 1938 -124 1972 -119
rect 2011 -124 2045 -119
rect 2084 -124 2118 -119
rect 2157 -124 2191 -119
rect 2230 -124 2264 -119
rect 2303 -124 2337 -119
rect 2376 -124 2410 -119
rect 2449 -124 2483 -119
rect 2522 -124 2556 -119
rect 2595 -124 2629 -119
rect 2668 -124 2702 -119
rect 1573 -153 1587 -124
rect 1587 -153 1607 -124
rect 1646 -153 1657 -124
rect 1657 -153 1680 -124
rect 1719 -153 1727 -124
rect 1727 -153 1753 -124
rect 1792 -153 1797 -124
rect 1797 -153 1826 -124
rect 1865 -153 1867 -124
rect 1867 -153 1899 -124
rect 1938 -153 1971 -124
rect 1971 -153 1972 -124
rect 2011 -153 2041 -124
rect 2041 -153 2045 -124
rect 2084 -153 2111 -124
rect 2111 -153 2118 -124
rect 2157 -153 2181 -124
rect 2181 -153 2191 -124
rect 2230 -153 2251 -124
rect 2251 -153 2264 -124
rect 2303 -153 2321 -124
rect 2321 -153 2337 -124
rect 2376 -153 2391 -124
rect 2391 -153 2410 -124
rect 2449 -153 2461 -124
rect 2461 -153 2483 -124
rect 2522 -153 2531 -124
rect 2531 -153 2556 -124
rect 2595 -153 2601 -124
rect 2601 -153 2629 -124
rect 2668 -153 2671 -124
rect 2671 -153 2702 -124
rect 2741 -153 2775 -119
rect 2814 -124 2848 -119
rect 2887 -124 2921 -119
rect 2960 -124 2994 -119
rect 3033 -124 3067 -119
rect 3106 -124 3140 -119
rect 3179 -124 3213 -119
rect 3252 -124 3286 -119
rect 3325 -124 3359 -119
rect 3398 -124 3432 -119
rect 3471 -124 3505 -119
rect 3544 -124 3578 -119
rect 3617 -124 3651 -119
rect 2814 -153 2847 -124
rect 2847 -153 2848 -124
rect 2887 -153 2917 -124
rect 2917 -153 2921 -124
rect 2960 -153 2987 -124
rect 2987 -153 2994 -124
rect 3033 -153 3057 -124
rect 3057 -153 3067 -124
rect 3106 -153 3127 -124
rect 3127 -153 3140 -124
rect 3179 -153 3197 -124
rect 3197 -153 3213 -124
rect 3252 -153 3267 -124
rect 3267 -153 3286 -124
rect 3325 -153 3337 -124
rect 3337 -153 3359 -124
rect 3398 -153 3407 -124
rect 3407 -153 3432 -124
rect 3471 -153 3477 -124
rect 3477 -153 3505 -124
rect 3544 -153 3547 -124
rect 3547 -153 3578 -124
rect 3617 -153 3651 -124
rect 3690 -153 3724 -119
rect 3763 -153 3797 -119
rect 3836 -153 3870 -119
rect 3909 -153 3943 -119
rect 3982 -153 4016 -119
rect 4055 -153 4089 -119
rect 4128 -153 4162 -119
rect 4201 -153 4235 -119
rect 4274 -153 4308 -119
rect 4347 -153 4381 -119
rect 4420 -153 4454 -119
rect 4493 -153 4527 -119
rect 4565 -153 4599 -119
rect 4637 -153 4671 -119
rect 4709 -153 4743 -119
rect 1573 -228 1587 -201
rect 1587 -228 1607 -201
rect 1646 -228 1657 -201
rect 1657 -228 1680 -201
rect 1719 -228 1727 -201
rect 1727 -228 1753 -201
rect 1792 -228 1797 -201
rect 1797 -228 1826 -201
rect 1865 -228 1867 -201
rect 1867 -228 1899 -201
rect 1938 -228 1971 -201
rect 1971 -228 1972 -201
rect 2011 -228 2041 -201
rect 2041 -228 2045 -201
rect 2084 -228 2111 -201
rect 2111 -228 2118 -201
rect 2157 -228 2181 -201
rect 2181 -228 2191 -201
rect 2230 -228 2251 -201
rect 2251 -228 2264 -201
rect 2303 -228 2321 -201
rect 2321 -228 2337 -201
rect 2376 -228 2391 -201
rect 2391 -228 2410 -201
rect 2449 -228 2461 -201
rect 2461 -228 2483 -201
rect 2522 -228 2531 -201
rect 2531 -228 2556 -201
rect 2595 -228 2601 -201
rect 2601 -228 2629 -201
rect 2668 -228 2671 -201
rect 2671 -228 2702 -201
rect 1573 -235 1607 -228
rect 1646 -235 1680 -228
rect 1719 -235 1753 -228
rect 1792 -235 1826 -228
rect 1865 -235 1899 -228
rect 1938 -235 1972 -228
rect 2011 -235 2045 -228
rect 2084 -235 2118 -228
rect 2157 -235 2191 -228
rect 2230 -235 2264 -228
rect 2303 -235 2337 -228
rect 2376 -235 2410 -228
rect 2449 -235 2483 -228
rect 2522 -235 2556 -228
rect 2595 -235 2629 -228
rect 2668 -235 2702 -228
rect 2741 -235 2775 -201
rect 2814 -228 2847 -201
rect 2847 -228 2848 -201
rect 2887 -228 2917 -201
rect 2917 -228 2921 -201
rect 2960 -228 2987 -201
rect 2987 -228 2994 -201
rect 3033 -228 3057 -201
rect 3057 -228 3067 -201
rect 3106 -228 3127 -201
rect 3127 -228 3140 -201
rect 3179 -228 3197 -201
rect 3197 -228 3213 -201
rect 3252 -228 3267 -201
rect 3267 -228 3286 -201
rect 3325 -228 3337 -201
rect 3337 -228 3359 -201
rect 3398 -228 3407 -201
rect 3407 -228 3432 -201
rect 3471 -228 3477 -201
rect 3477 -228 3505 -201
rect 3544 -228 3547 -201
rect 3547 -228 3578 -201
rect 3617 -228 3651 -201
rect 2814 -235 2848 -228
rect 2887 -235 2921 -228
rect 2960 -235 2994 -228
rect 3033 -235 3067 -228
rect 3106 -235 3140 -228
rect 3179 -235 3213 -228
rect 3252 -235 3286 -228
rect 3325 -235 3359 -228
rect 3398 -235 3432 -228
rect 3471 -235 3505 -228
rect 3544 -235 3578 -228
rect 3617 -235 3651 -228
rect 3690 -235 3724 -201
rect 3763 -235 3797 -201
rect 3836 -235 3870 -201
rect 3909 -235 3943 -201
rect 3982 -235 4016 -201
rect 4055 -235 4089 -201
rect 4128 -235 4162 -201
rect 4201 -235 4235 -201
rect 4274 -235 4308 -201
rect 4347 -235 4381 -201
rect 4420 -235 4454 -201
rect 4493 -235 4527 -201
rect 4565 -235 4599 -201
rect 4637 -235 4671 -201
rect 4709 -235 4743 -201
rect 1480 -946 1514 -912
rect 1556 -928 1587 -912
rect 1587 -928 1590 -912
rect 1632 -928 1657 -912
rect 1657 -928 1666 -912
rect 1707 -928 1727 -912
rect 1727 -928 1741 -912
rect 1782 -928 1797 -912
rect 1797 -928 1816 -912
rect 1857 -928 1867 -912
rect 1867 -928 1891 -912
rect 1932 -928 1937 -912
rect 1937 -928 1966 -912
rect 2007 -928 2041 -912
rect 2082 -928 2111 -912
rect 2111 -928 2116 -912
rect 2157 -928 2181 -912
rect 2181 -928 2191 -912
rect 2232 -928 2251 -912
rect 2251 -928 2266 -912
rect 2307 -928 2321 -912
rect 2321 -928 2341 -912
rect 2382 -928 2391 -912
rect 2391 -928 2416 -912
rect 2457 -928 2461 -912
rect 2461 -928 2491 -912
rect 1556 -946 1590 -928
rect 1632 -946 1666 -928
rect 1707 -946 1741 -928
rect 1782 -946 1816 -928
rect 1857 -946 1891 -928
rect 1932 -946 1966 -928
rect 2007 -946 2041 -928
rect 2082 -946 2116 -928
rect 2157 -946 2191 -928
rect 2232 -946 2266 -928
rect 2307 -946 2341 -928
rect 2382 -946 2416 -928
rect 2457 -946 2491 -928
rect 2532 -946 2566 -912
rect 2607 -928 2637 -912
rect 2637 -928 2641 -912
rect 2682 -928 2707 -912
rect 2707 -928 2716 -912
rect 2757 -928 2777 -912
rect 2777 -928 2791 -912
rect 2832 -928 2847 -912
rect 2847 -928 2866 -912
rect 2907 -928 2917 -912
rect 2917 -928 2941 -912
rect 2982 -928 2987 -912
rect 2987 -928 3016 -912
rect 3057 -928 3091 -912
rect 3132 -928 3161 -912
rect 3161 -928 3166 -912
rect 3207 -928 3231 -912
rect 3231 -928 3241 -912
rect 2607 -946 2641 -928
rect 2682 -946 2716 -928
rect 2757 -946 2791 -928
rect 2832 -946 2866 -928
rect 2907 -946 2941 -928
rect 2982 -946 3016 -928
rect 3057 -946 3091 -928
rect 3132 -946 3166 -928
rect 3207 -946 3241 -928
<< metal1 >>
rect 10582 2510 10588 2562
rect 10640 2510 10660 2562
rect 10712 2510 10732 2562
rect 10784 2510 10803 2562
rect 10855 2510 10861 2562
rect 10582 2490 10861 2510
rect 10582 2438 10588 2490
rect 10640 2438 10660 2490
rect 10712 2438 10732 2490
rect 10784 2438 10803 2490
rect 10855 2438 10861 2490
rect -179 2033 -139 2235
rect 10582 2234 10861 2235
rect 10582 2182 10588 2234
rect 10640 2182 10660 2234
rect 10712 2182 10732 2234
rect 10784 2182 10803 2234
rect 10855 2182 10861 2234
rect 10582 2160 10861 2182
rect 10582 2108 10588 2160
rect 10640 2108 10660 2160
rect 10712 2108 10732 2160
rect 10784 2108 10803 2160
rect 10855 2108 10861 2160
rect 10582 2086 10861 2108
rect 10582 2034 10588 2086
rect 10640 2034 10660 2086
rect 10712 2034 10732 2086
rect 10784 2034 10803 2086
rect 10855 2034 10861 2086
rect 10582 2033 10861 2034
rect 12524 2033 12564 2235
rect 54 1875 94 2005
rect 104 1998 220 2004
rect 104 1876 220 1882
rect 2570 1999 3714 2005
rect 2570 1965 2582 1999
rect 2616 1965 2655 1999
rect 2689 1965 2728 1999
rect 2762 1965 2801 1999
rect 2835 1965 2874 1999
rect 2908 1965 2947 1999
rect 2981 1965 3020 1999
rect 3054 1965 3092 1999
rect 3126 1965 3164 1999
rect 3198 1965 3236 1999
rect 3270 1965 3308 1999
rect 3342 1965 3380 1999
rect 3414 1965 3452 1999
rect 3486 1965 3524 1999
rect 3558 1965 3596 1999
rect 3630 1965 3668 1999
rect 3702 1965 3714 1999
rect 2570 1915 3714 1965
rect 2570 1881 2582 1915
rect 2616 1881 2655 1915
rect 2689 1881 2728 1915
rect 2762 1881 2801 1915
rect 2835 1881 2874 1915
rect 2908 1881 2947 1915
rect 2981 1881 3020 1915
rect 3054 1881 3092 1915
rect 3126 1881 3164 1915
rect 3198 1881 3236 1915
rect 3270 1881 3308 1915
rect 3342 1881 3380 1915
rect 3414 1881 3452 1915
rect 3486 1881 3524 1915
rect 3558 1881 3596 1915
rect 3630 1881 3668 1915
rect 3702 1881 3714 1915
rect 2570 1875 3714 1881
rect 3732 1953 3738 2005
rect 3790 1953 3809 2005
rect 3861 1953 3880 2005
rect 3932 1953 3950 2005
rect 4002 1953 4020 2005
rect 4072 1953 4090 2005
rect 4142 1953 4160 2005
rect 4212 1953 4230 2005
rect 4282 1953 4288 2005
rect 3732 1927 4288 1953
rect 3732 1875 3738 1927
rect 3790 1875 3809 1927
rect 3861 1875 3880 1927
rect 3932 1875 3950 1927
rect 4002 1875 4020 1927
rect 4072 1875 4090 1927
rect 4142 1875 4160 1927
rect 4212 1875 4230 1927
rect 4282 1875 4288 1927
rect 7927 1953 7933 2005
rect 7985 1953 8037 2005
rect 8089 1953 8141 2005
rect 8193 1953 8245 2005
rect 8297 1953 8348 2005
rect 8400 1953 8451 2005
rect 8503 1953 8509 2005
rect 7927 1927 8509 1953
rect 7927 1875 7933 1927
rect 7985 1875 8037 1927
rect 8089 1875 8141 1927
rect 8193 1875 8245 1927
rect 8297 1875 8348 1927
rect 8400 1875 8451 1927
rect 8503 1875 8509 1927
rect 12433 1875 12473 2005
rect 2073 1792 4702 1797
rect 7816 1795 7866 1847
rect 2073 1740 2084 1792
rect 2136 1740 2148 1792
rect 2200 1740 4580 1792
rect 4632 1740 4644 1792
rect 4696 1740 4702 1792
rect 2073 1737 4702 1740
rect 7493 1715 7545 1767
rect 476 1583 6798 1589
rect 476 1549 488 1583
rect 522 1549 560 1583
rect 594 1549 6746 1583
rect 476 1543 6746 1549
tri 6721 1518 6746 1543 ne
rect 6746 1519 6798 1531
rect 6226 1443 6232 1495
rect 6284 1443 6296 1495
rect 6348 1443 6368 1495
rect 6746 1461 6798 1467
tri 6240 1415 6268 1443 ne
rect 6268 1287 6368 1443
tri 6726 1287 6750 1311 se
rect 6750 1287 11121 1311
rect 6267 1276 11121 1287
tri 11121 1276 11156 1311 sw
rect 6267 1268 11156 1276
rect 6267 1235 6735 1268
tri 6735 1235 6768 1268 nw
tri 11107 1235 11140 1268 ne
rect 11140 1235 11156 1268
tri 11140 1219 11156 1235 ne
tri 11156 1219 11213 1276 sw
tri 11156 1213 11162 1219 ne
rect 11162 1213 12335 1219
tri 11162 1207 11168 1213 ne
rect 11168 1207 11785 1213
rect 5785 1201 6378 1207
rect 5785 1167 5797 1201
rect 5831 1167 5869 1201
rect 5903 1167 6378 1201
rect 5785 1161 6378 1167
tri 6358 1152 6367 1161 ne
rect 6367 1152 6378 1161
tri 6378 1152 6433 1207 sw
tri 11168 1176 11199 1207 ne
rect 11199 1176 11785 1207
tri 11748 1152 11772 1176 ne
rect 11772 1152 11785 1176
tri 6367 1141 6378 1152 ne
rect 6378 1141 6433 1152
tri 6378 1107 6412 1141 ne
rect 6412 1107 6433 1141
tri 6433 1107 6478 1152 sw
tri 11772 1151 11773 1152 ne
rect 11773 1107 11785 1152
rect 12323 1107 12335 1213
tri 6412 1086 6433 1107 ne
rect 6433 1086 6478 1107
tri 6478 1086 6499 1107 sw
rect 11773 1101 12335 1107
rect -179 884 -96 1086
rect 104 1080 220 1086
rect 156 1028 168 1080
rect 3080 1080 3226 1086
rect 104 1008 220 1028
rect 156 956 168 1008
rect 104 936 220 956
rect 156 884 168 936
rect 862 1052 908 1064
rect 862 1018 868 1052
rect 902 1018 908 1052
rect 862 980 908 1018
rect 862 946 868 980
rect 902 946 908 980
rect 862 934 908 946
rect 3132 1028 3174 1080
rect 3080 1011 3226 1028
rect 3132 959 3174 1011
rect 3080 942 3226 959
rect 3132 890 3174 942
rect 3080 884 3226 890
rect 3732 1034 3738 1086
rect 3790 1034 3809 1086
rect 3861 1034 3880 1086
rect 3932 1034 3950 1086
rect 4002 1034 4020 1086
rect 4072 1034 4090 1086
rect 4142 1034 4160 1086
rect 4212 1034 4230 1086
rect 4282 1034 4288 1086
tri 6433 1074 6445 1086 ne
rect 6445 1074 7090 1086
tri 6445 1058 6461 1074 ne
rect 6461 1058 7050 1074
tri 7019 1052 7025 1058 ne
rect 7025 1052 7050 1058
rect 3732 1011 4288 1034
rect 3732 959 3738 1011
rect 3790 959 3809 1011
rect 3861 959 3880 1011
rect 3932 959 3950 1011
rect 4002 959 4020 1011
rect 4072 959 4090 1011
rect 4142 959 4160 1011
rect 4212 959 4230 1011
rect 4282 959 4288 1011
rect 3732 936 4288 959
rect 3732 884 3738 936
rect 3790 884 3809 936
rect 3861 884 3880 936
rect 3932 884 3950 936
rect 4002 884 4020 936
rect 4072 884 4090 936
rect 4142 884 4160 936
rect 4212 884 4230 936
rect 4282 884 4288 936
rect 5388 1040 5434 1052
tri 7025 1040 7037 1052 ne
rect 7037 1040 7050 1052
rect 7084 1040 7090 1074
rect 5388 1006 5394 1040
rect 5428 1006 5434 1040
tri 7037 1033 7044 1040 ne
rect 5388 968 5434 1006
rect 5388 934 5394 968
rect 5428 934 5434 968
rect 5388 922 5434 934
rect 6633 1024 6798 1030
rect 6633 972 6746 1024
rect 6633 960 6798 972
rect 6633 908 6746 960
rect 7044 1002 7090 1040
rect 7044 968 7050 1002
rect 7084 968 7090 1002
rect 7044 956 7090 968
rect 6633 900 6798 908
tri 5883 884 5884 885 ne
rect 5884 884 6049 885
rect 104 865 220 884
rect 156 813 168 865
tri 5884 850 5918 884 ne
rect 5918 850 6049 884
tri 6049 850 6083 884 nw
tri 5918 845 5923 850 ne
rect 5923 845 6049 850
tri 5923 815 5953 845 ne
rect 5953 815 6049 845
rect 104 794 220 813
tri 5953 802 5966 815 ne
rect 156 742 168 794
rect 104 736 220 742
rect 5966 784 6049 815
tri 6049 784 6080 815 sw
rect 7927 793 7933 845
rect 7985 793 8016 845
rect 8068 793 8099 845
rect 8151 793 8181 845
rect 8233 793 8263 845
rect 8315 793 8345 845
rect 8397 793 8403 845
rect 5966 740 6156 784
tri 6156 740 6200 784 sw
rect 7927 770 8403 793
rect 5966 697 6224 740
rect 7927 718 7933 770
rect 7985 718 8016 770
rect 8068 718 8099 770
rect 8151 718 8181 770
rect 8233 718 8263 770
rect 8315 718 8345 770
rect 8397 718 8403 770
tri 6224 697 6243 716 sw
rect 5966 692 6243 697
rect 7927 695 8403 718
rect 5212 630 5535 636
rect 5212 624 5483 630
rect 5212 590 5218 624
rect 5252 590 5483 624
rect 5212 578 5483 590
rect 5212 564 5535 578
rect 5212 552 5483 564
rect 5212 518 5218 552
rect 5252 518 5483 552
rect 5212 512 5483 518
rect 5212 506 5535 512
rect 5684 630 5736 636
rect 5684 564 5736 578
rect 3065 239 3231 441
rect 5367 239 5434 441
rect 5591 369 5637 478
rect 5684 392 5736 512
rect 5966 478 6224 692
rect 7927 643 7933 695
rect 7985 643 8016 695
rect 8068 643 8099 695
rect 8151 643 8181 695
rect 8233 643 8263 695
rect 8315 643 8345 695
rect 8397 643 8403 695
tri 5684 377 5699 392 ne
rect 5699 377 5736 392
tri 5637 369 5645 377 sw
tri 5699 369 5707 377 ne
rect 5707 369 5736 377
tri 5736 369 5781 414 sw
rect 5591 357 5645 369
tri 5645 357 5657 369 sw
tri 5707 357 5719 369 ne
rect 5719 357 6804 369
tri 5591 340 5608 357 ne
rect 5608 348 5657 357
tri 5657 348 5666 357 sw
rect 5608 340 5666 348
tri 5719 340 5736 357 ne
rect 5736 340 6804 357
tri 5608 334 5614 340 ne
rect 738 211 5499 239
rect 5614 223 5666 340
tri 5736 317 5759 340 ne
rect 5759 317 6804 340
rect 5367 93 5434 211
rect 1771 -15 2052 -9
rect 1771 -49 1783 -15
rect 1817 -49 1855 -15
rect 1889 -49 2052 -15
rect 1771 -55 2052 -49
tri 2040 -59 2044 -55 ne
rect 2044 -59 2052 -55
tri 2044 -61 2046 -59 ne
rect 2046 -61 2052 -59
rect 2104 -61 2116 -9
rect 2168 -61 2174 -9
tri 2995 -41 3018 -18 se
rect 3018 -21 3024 31
rect 3076 -21 3093 31
rect 3145 -7 3161 31
rect 3213 -21 3229 31
rect 3281 -21 3287 31
rect 3018 -41 3030 -21
rect 3064 -41 3136 -21
rect 3170 -41 3241 -21
rect 3275 -25 3287 -21
tri 3287 -25 3297 -15 sw
rect 3275 -41 3297 -25
tri 2977 -59 2995 -41 se
rect 2995 -49 3297 -41
tri 3297 -49 3321 -25 sw
rect 4571 -49 4580 3
rect 4632 -49 4644 3
rect 4696 -49 4702 3
rect 2995 -59 3321 -49
tri 3321 -59 3331 -49 sw
rect 4571 -59 4583 -49
rect 4617 -59 4655 -49
rect 4689 -59 4702 -49
tri 2975 -61 2977 -59 se
rect 2977 -61 3331 -59
tri 2923 -113 2975 -61 se
rect 2975 -63 3331 -61
rect 2975 -113 3024 -63
rect 1561 -115 3024 -113
rect 3076 -115 3093 -63
rect 3145 -115 3161 -63
rect 3213 -115 3229 -63
rect 3281 -65 3331 -63
tri 3331 -65 3337 -59 sw
rect 4571 -65 4702 -59
rect 3281 -113 3337 -65
tri 3337 -113 3385 -65 sw
rect 3281 -115 4755 -113
rect 1561 -119 4755 -115
rect 1561 -153 1573 -119
rect 1607 -153 1646 -119
rect 1680 -153 1719 -119
rect 1753 -153 1792 -119
rect 1826 -153 1865 -119
rect 1899 -153 1938 -119
rect 1972 -153 2011 -119
rect 2045 -153 2084 -119
rect 2118 -153 2157 -119
rect 2191 -153 2230 -119
rect 2264 -153 2303 -119
rect 2337 -153 2376 -119
rect 2410 -153 2449 -119
rect 2483 -153 2522 -119
rect 2556 -153 2595 -119
rect 2629 -153 2668 -119
rect 2702 -153 2741 -119
rect 2775 -153 2814 -119
rect 2848 -153 2887 -119
rect 2921 -153 2960 -119
rect 2994 -153 3033 -119
rect 3067 -153 3106 -119
rect 3140 -153 3179 -119
rect 3213 -153 3252 -119
rect 3286 -153 3325 -119
rect 3359 -153 3398 -119
rect 3432 -153 3471 -119
rect 3505 -153 3544 -119
rect 3578 -153 3617 -119
rect 3651 -153 3690 -119
rect 3724 -153 3763 -119
rect 3797 -153 3836 -119
rect 3870 -153 3909 -119
rect 3943 -153 3982 -119
rect 4016 -153 4055 -119
rect 4089 -153 4128 -119
rect 4162 -153 4201 -119
rect 4235 -153 4274 -119
rect 4308 -153 4347 -119
rect 4381 -153 4420 -119
rect 4454 -153 4493 -119
rect 4527 -153 4565 -119
rect 4599 -153 4637 -119
rect 4671 -153 4709 -119
rect 4743 -153 4755 -119
rect 1561 -201 4755 -153
rect 1561 -235 1573 -201
rect 1607 -235 1646 -201
rect 1680 -235 1719 -201
rect 1753 -235 1792 -201
rect 1826 -235 1865 -201
rect 1899 -235 1938 -201
rect 1972 -235 2011 -201
rect 2045 -235 2084 -201
rect 2118 -235 2157 -201
rect 2191 -235 2230 -201
rect 2264 -235 2303 -201
rect 2337 -235 2376 -201
rect 2410 -235 2449 -201
rect 2483 -235 2522 -201
rect 2556 -235 2595 -201
rect 2629 -235 2668 -201
rect 2702 -235 2741 -201
rect 2775 -235 2814 -201
rect 2848 -235 2887 -201
rect 2921 -235 2960 -201
rect 2994 -235 3033 -201
rect 3067 -235 3106 -201
rect 3140 -235 3179 -201
rect 3213 -235 3252 -201
rect 3286 -235 3325 -201
rect 3359 -235 3398 -201
rect 3432 -235 3471 -201
rect 3505 -235 3544 -201
rect 3578 -235 3617 -201
rect 3651 -235 3690 -201
rect 3724 -235 3763 -201
rect 3797 -235 3836 -201
rect 3870 -235 3909 -201
rect 3943 -235 3982 -201
rect 4016 -235 4055 -201
rect 4089 -235 4128 -201
rect 4162 -235 4201 -201
rect 4235 -235 4274 -201
rect 4308 -235 4347 -201
rect 4381 -235 4420 -201
rect 4454 -235 4493 -201
rect 4527 -235 4565 -201
rect 4599 -235 4637 -201
rect 4671 -235 4709 -201
rect 4743 -235 4755 -201
rect 1561 -241 4755 -235
tri 1788 -906 1791 -903 se
rect 1791 -906 1797 -903
rect 1468 -912 1797 -906
rect 1849 -912 1865 -903
rect 1917 -912 1933 -903
rect 1468 -946 1480 -912
rect 1514 -946 1556 -912
rect 1590 -946 1632 -912
rect 1666 -946 1707 -912
rect 1741 -946 1782 -912
rect 1849 -946 1857 -912
rect 1917 -946 1932 -912
rect 1468 -952 1797 -946
tri 1788 -955 1791 -952 ne
rect 1791 -955 1797 -952
rect 1849 -955 1865 -946
rect 1917 -955 1933 -946
rect 1985 -955 2001 -903
rect 2053 -955 2069 -903
rect 2121 -955 2137 -903
rect 2189 -912 2205 -903
rect 2257 -912 2273 -903
rect 2325 -906 2331 -903
tri 2331 -906 2334 -903 sw
rect 2325 -912 3253 -906
rect 2191 -946 2205 -912
rect 2266 -946 2273 -912
rect 2341 -946 2382 -912
rect 2416 -946 2457 -912
rect 2491 -946 2532 -912
rect 2566 -946 2607 -912
rect 2641 -946 2682 -912
rect 2716 -946 2757 -912
rect 2791 -946 2832 -912
rect 2866 -946 2907 -912
rect 2941 -946 2982 -912
rect 3016 -946 3057 -912
rect 3091 -946 3132 -912
rect 3166 -946 3207 -912
rect 3241 -946 3253 -912
rect 2189 -955 2205 -946
rect 2257 -955 2273 -946
rect 2325 -952 3253 -946
rect 2325 -955 2331 -952
tri 2331 -955 2334 -952 nw
<< via1 >>
rect 10588 2510 10640 2562
rect 10660 2510 10712 2562
rect 10732 2510 10784 2562
rect 10803 2510 10855 2562
rect 10588 2438 10640 2490
rect 10660 2438 10712 2490
rect 10732 2438 10784 2490
rect 10803 2438 10855 2490
rect 10588 2182 10640 2234
rect 10660 2182 10712 2234
rect 10732 2182 10784 2234
rect 10803 2182 10855 2234
rect 10588 2108 10640 2160
rect 10660 2108 10712 2160
rect 10732 2108 10784 2160
rect 10803 2108 10855 2160
rect 10588 2034 10640 2086
rect 10660 2034 10712 2086
rect 10732 2034 10784 2086
rect 10803 2034 10855 2086
rect 104 1882 220 1998
rect 3738 1953 3790 2005
rect 3809 1953 3861 2005
rect 3880 1953 3932 2005
rect 3950 1953 4002 2005
rect 4020 1953 4072 2005
rect 4090 1953 4142 2005
rect 4160 1953 4212 2005
rect 4230 1953 4282 2005
rect 3738 1875 3790 1927
rect 3809 1875 3861 1927
rect 3880 1875 3932 1927
rect 3950 1875 4002 1927
rect 4020 1875 4072 1927
rect 4090 1875 4142 1927
rect 4160 1875 4212 1927
rect 4230 1875 4282 1927
rect 7933 1953 7985 2005
rect 8037 1953 8089 2005
rect 8141 1953 8193 2005
rect 8245 1953 8297 2005
rect 8348 1953 8400 2005
rect 8451 1953 8503 2005
rect 7933 1875 7985 1927
rect 8037 1875 8089 1927
rect 8141 1875 8193 1927
rect 8245 1875 8297 1927
rect 8348 1875 8400 1927
rect 8451 1875 8503 1927
rect 2084 1740 2136 1792
rect 2148 1740 2200 1792
rect 4580 1740 4632 1792
rect 4644 1740 4696 1792
rect 6746 1531 6798 1583
rect 6232 1443 6284 1495
rect 6296 1443 6348 1495
rect 6746 1467 6798 1519
rect 104 1028 156 1080
rect 168 1028 220 1080
rect 104 956 156 1008
rect 168 956 220 1008
rect 104 884 156 936
rect 168 884 220 936
rect 3080 1028 3132 1080
rect 3174 1028 3226 1080
rect 3080 959 3132 1011
rect 3174 959 3226 1011
rect 3080 890 3132 942
rect 3174 890 3226 942
rect 3738 1034 3790 1086
rect 3809 1034 3861 1086
rect 3880 1034 3932 1086
rect 3950 1034 4002 1086
rect 4020 1034 4072 1086
rect 4090 1034 4142 1086
rect 4160 1034 4212 1086
rect 4230 1034 4282 1086
rect 3738 959 3790 1011
rect 3809 959 3861 1011
rect 3880 959 3932 1011
rect 3950 959 4002 1011
rect 4020 959 4072 1011
rect 4090 959 4142 1011
rect 4160 959 4212 1011
rect 4230 959 4282 1011
rect 3738 884 3790 936
rect 3809 884 3861 936
rect 3880 884 3932 936
rect 3950 884 4002 936
rect 4020 884 4072 936
rect 4090 884 4142 936
rect 4160 884 4212 936
rect 4230 884 4282 936
rect 6746 972 6798 1024
rect 6746 908 6798 960
rect 104 813 156 865
rect 168 813 220 865
rect 104 742 156 794
rect 168 742 220 794
rect 7933 793 7985 845
rect 8016 793 8068 845
rect 8099 793 8151 845
rect 8181 793 8233 845
rect 8263 793 8315 845
rect 8345 793 8397 845
rect 7933 718 7985 770
rect 8016 718 8068 770
rect 8099 718 8151 770
rect 8181 718 8233 770
rect 8263 718 8315 770
rect 8345 718 8397 770
rect 5483 578 5535 630
rect 5483 512 5535 564
rect 5684 578 5736 630
rect 5684 512 5736 564
rect 7933 643 7985 695
rect 8016 643 8068 695
rect 8099 643 8151 695
rect 8181 643 8233 695
rect 8263 643 8315 695
rect 8345 643 8397 695
rect 2052 -61 2104 -9
rect 2116 -61 2168 -9
rect 3024 -7 3076 31
rect 3024 -21 3030 -7
rect 3030 -21 3064 -7
rect 3064 -21 3076 -7
rect 3093 -7 3145 31
rect 3161 -7 3213 31
rect 3093 -21 3136 -7
rect 3136 -21 3145 -7
rect 3161 -21 3170 -7
rect 3170 -21 3213 -7
rect 3229 -7 3281 31
rect 3229 -21 3241 -7
rect 3241 -21 3275 -7
rect 3275 -21 3281 -7
rect 4580 -25 4632 3
rect 4580 -49 4583 -25
rect 4583 -49 4617 -25
rect 4617 -49 4632 -25
rect 4644 -25 4696 3
rect 4644 -49 4655 -25
rect 4655 -49 4689 -25
rect 4689 -49 4696 -25
rect 3024 -115 3076 -63
rect 3093 -115 3145 -63
rect 3161 -115 3213 -63
rect 3229 -115 3281 -63
rect 1797 -912 1849 -903
rect 1865 -912 1917 -903
rect 1933 -912 1985 -903
rect 1797 -946 1816 -912
rect 1816 -946 1849 -912
rect 1865 -946 1891 -912
rect 1891 -946 1917 -912
rect 1933 -946 1966 -912
rect 1966 -946 1985 -912
rect 1797 -955 1849 -946
rect 1865 -955 1917 -946
rect 1933 -955 1985 -946
rect 2001 -912 2053 -903
rect 2001 -946 2007 -912
rect 2007 -946 2041 -912
rect 2041 -946 2053 -912
rect 2001 -955 2053 -946
rect 2069 -912 2121 -903
rect 2069 -946 2082 -912
rect 2082 -946 2116 -912
rect 2116 -946 2121 -912
rect 2069 -955 2121 -946
rect 2137 -912 2189 -903
rect 2205 -912 2257 -903
rect 2273 -912 2325 -903
rect 2137 -946 2157 -912
rect 2157 -946 2189 -912
rect 2205 -946 2232 -912
rect 2232 -946 2257 -912
rect 2273 -946 2307 -912
rect 2307 -946 2325 -912
rect 2137 -955 2189 -946
rect 2205 -955 2257 -946
rect 2273 -955 2325 -946
<< metal2 >>
rect 10582 2510 10588 2562
rect 10640 2510 10660 2562
rect 10712 2510 10732 2562
rect 10784 2510 10803 2562
rect 10855 2510 10861 2562
rect 10582 2490 10861 2510
rect 10582 2438 10588 2490
rect 10640 2438 10660 2490
rect 10712 2438 10732 2490
rect 10784 2438 10803 2490
rect 10855 2438 10861 2490
rect 10582 2234 10861 2438
rect 10582 2182 10588 2234
rect 10640 2182 10660 2234
rect 10712 2182 10732 2234
rect 10784 2182 10803 2234
rect 10855 2182 10861 2234
rect 10582 2160 10861 2182
rect 10582 2108 10588 2160
rect 10640 2108 10660 2160
rect 10712 2108 10732 2160
rect 10784 2108 10803 2160
rect 10855 2108 10861 2160
rect 10582 2086 10861 2108
rect 10582 2034 10588 2086
rect 10640 2034 10660 2086
rect 10712 2034 10732 2086
rect 10784 2034 10803 2086
rect 10855 2034 10861 2086
rect 10582 2033 10861 2034
rect 104 1998 220 2004
rect 104 1080 220 1882
rect 3732 1953 3738 2005
rect 3790 1953 3809 2005
rect 3861 1953 3880 2005
rect 3932 1953 3950 2005
rect 4002 1953 4020 2005
rect 4072 1953 4090 2005
rect 4142 1953 4160 2005
rect 4212 1953 4230 2005
rect 4282 1953 4288 2005
rect 3732 1927 4288 1953
rect 3732 1875 3738 1927
rect 3790 1875 3809 1927
rect 3861 1875 3880 1927
rect 3932 1875 3950 1927
rect 4002 1875 4020 1927
rect 4072 1875 4090 1927
rect 4142 1875 4160 1927
rect 4212 1875 4230 1927
rect 4282 1875 4288 1927
rect 7927 1953 7933 2005
rect 7985 1968 8037 2005
rect 8089 1968 8141 2005
rect 8193 1968 8245 2005
rect 8297 1968 8348 2005
rect 8400 1968 8451 2005
rect 7992 1953 8037 1968
rect 7927 1927 7936 1953
rect 7992 1927 8038 1953
rect 7927 1875 7933 1927
rect 7992 1912 8037 1927
rect 8094 1912 8140 1968
rect 8196 1912 8242 1968
rect 8298 1912 8343 1968
rect 8400 1953 8444 1968
rect 8503 1953 8509 2005
rect 8399 1927 8444 1953
rect 8500 1927 8509 1953
rect 8400 1912 8444 1927
rect 7985 1875 8037 1912
rect 8089 1875 8141 1912
rect 8193 1875 8245 1912
rect 8297 1875 8348 1912
rect 8400 1875 8451 1912
rect 8503 1875 8509 1927
tri 1848 1740 1900 1792 se
rect 1900 1740 2084 1792
rect 2136 1740 2148 1792
rect 2200 1740 2206 1792
tri 1813 1705 1848 1740 se
rect 1848 1705 1887 1740
tri 1887 1705 1922 1740 nw
tri 1739 1631 1813 1705 se
tri 1813 1631 1887 1705 nw
tri 1691 1583 1739 1631 se
rect 1739 1583 1765 1631
tri 1765 1583 1813 1631 nw
tri 1665 1557 1691 1583 se
rect 1691 1557 1739 1583
tri 1739 1557 1765 1583 nw
tri 1639 1531 1665 1557 se
rect 1665 1531 1713 1557
tri 1713 1531 1739 1557 nw
tri 1627 1519 1639 1531 se
rect 1639 1519 1701 1531
tri 1701 1519 1713 1531 nw
tri 1603 1495 1627 1519 se
rect 1627 1495 1677 1519
tri 1677 1495 1701 1519 nw
tri 1591 1483 1603 1495 se
rect 1603 1483 1665 1495
tri 1665 1483 1677 1495 nw
tri 1551 1443 1591 1483 se
rect 1591 1443 1625 1483
tri 1625 1443 1665 1483 nw
tri 1517 1409 1551 1443 se
rect 1551 1409 1591 1443
tri 1591 1409 1625 1443 nw
rect 156 1028 168 1080
rect 104 1008 220 1028
rect 156 956 168 1008
rect 104 936 220 956
rect 156 884 168 936
rect 104 865 220 884
rect 156 813 168 865
tri 1465 1357 1517 1409 se
rect 1465 855 1517 1357
tri 1517 1335 1591 1409 nw
rect 3080 1080 3226 1087
rect 3132 1028 3174 1080
rect 3080 1011 3226 1028
rect 3132 959 3174 1011
rect 3080 942 3226 959
rect 3132 890 3174 942
tri 1465 854 1466 855 ne
rect 1466 854 1517 855
tri 1517 854 1540 877 sw
tri 1466 845 1475 854 ne
rect 1475 845 1540 854
tri 1540 845 1549 854 sw
rect 104 794 220 813
tri 1475 803 1517 845 ne
rect 1517 803 1549 845
rect 156 742 168 794
tri 1517 793 1527 803 ne
rect 1527 793 1549 803
tri 1549 793 1601 845 sw
tri 1527 780 1540 793 ne
rect 1540 780 1601 793
tri 1601 780 1614 793 sw
tri 1540 770 1550 780 ne
rect 1550 770 1614 780
tri 1614 770 1624 780 sw
rect 104 736 220 742
tri 1550 736 1584 770 ne
rect 1584 736 1624 770
tri 1584 718 1602 736 ne
rect 1602 718 1624 736
tri 1624 718 1676 770 sw
tri 1602 706 1614 718 ne
rect 1614 706 1676 718
tri 1676 706 1688 718 sw
tri 1614 695 1625 706 ne
rect 1625 695 2056 706
tri 2056 695 2067 706 sw
tri 1625 662 1658 695 ne
rect 1658 662 2067 695
tri 2067 662 2100 695 sw
tri 1658 654 1666 662 ne
rect 1666 654 2100 662
tri 2034 643 2045 654 ne
rect 2045 643 2100 654
tri 2100 643 2119 662 sw
tri 2045 630 2058 643 ne
rect 2058 630 2119 643
tri 2119 630 2132 643 sw
tri 2058 588 2100 630 ne
rect 2100 588 2132 630
tri 2132 588 2174 630 sw
tri 2100 578 2110 588 ne
rect 2110 578 2174 588
tri 2110 569 2119 578 ne
tri 2086 31 2119 64 se
rect 2119 31 2174 578
tri 3079 92 3080 93 se
rect 3080 92 3226 890
rect 3732 1086 4288 1875
rect 4571 1740 4580 1792
rect 4632 1740 4644 1792
rect 4696 1740 4702 1792
tri 4571 1721 4590 1740 ne
rect 3732 1034 3738 1086
rect 3790 1034 3809 1086
rect 3861 1034 3880 1086
rect 3932 1034 3950 1086
rect 4002 1034 4020 1086
rect 4072 1034 4090 1086
rect 4142 1034 4160 1086
rect 4212 1034 4230 1086
rect 4282 1034 4288 1086
rect 3732 1011 4288 1034
rect 3732 959 3738 1011
rect 3790 959 3809 1011
rect 3861 959 3880 1011
rect 3932 959 3950 1011
rect 4002 959 4020 1011
rect 4072 959 4090 1011
rect 4142 959 4160 1011
rect 4212 959 4230 1011
rect 4282 959 4288 1011
rect 3732 936 4288 959
rect 3732 884 3738 936
rect 3790 884 3809 936
rect 3861 884 3880 936
rect 3932 884 3950 936
rect 4002 884 4020 936
rect 4072 884 4090 936
rect 4142 884 4160 936
rect 4212 884 4230 936
rect 4282 884 4288 936
tri 3052 65 3079 92 se
rect 3079 65 3226 92
tri 2046 -9 2086 31 se
rect 2086 -9 2174 31
rect 2887 19 2933 65
tri 3018 31 3052 65 se
rect 3052 31 3226 65
tri 3226 31 3287 92 sw
rect 2046 -61 2052 -9
rect 2104 -61 2116 -9
rect 2168 -61 2174 -9
rect 3018 -21 3024 31
rect 3076 -21 3093 31
rect 3145 -21 3161 31
rect 3213 -21 3229 31
rect 3281 -21 3287 31
rect 3360 19 3411 49
tri 4587 19 4590 22 se
rect 4590 19 4668 1740
tri 4668 1706 4702 1740 nw
rect 6746 1583 6798 1589
rect 6746 1519 6798 1531
rect 6226 1443 6232 1495
rect 6284 1443 6296 1495
rect 6348 1443 6354 1495
rect 6746 1024 6798 1467
rect 6746 960 6798 972
rect 6746 902 6798 908
rect 7927 793 7933 845
rect 7985 840 8016 845
rect 8068 840 8099 845
rect 8151 840 8181 845
rect 8233 840 8263 845
rect 8315 840 8345 845
rect 7992 793 8016 840
rect 8091 793 8099 840
rect 8315 793 8332 840
rect 8397 793 8403 845
rect 7927 784 7936 793
rect 7992 784 8035 793
rect 8091 784 8134 793
rect 8190 784 8233 793
rect 8289 784 8332 793
rect 8388 784 8403 793
rect 7927 770 8403 784
rect 7927 718 7933 770
rect 7985 760 8016 770
rect 8068 760 8099 770
rect 8151 760 8181 770
rect 8233 760 8263 770
rect 8315 760 8345 770
rect 7992 718 8016 760
rect 8091 718 8099 760
rect 8315 718 8332 760
rect 8397 718 8403 770
rect 7927 704 7936 718
rect 7992 704 8035 718
rect 8091 704 8134 718
rect 8190 704 8233 718
rect 8289 704 8332 718
rect 8388 704 8403 718
rect 7927 695 8403 704
rect 7927 643 7933 695
rect 7985 643 8016 695
rect 8068 643 8099 695
rect 8151 643 8181 695
rect 8233 643 8263 695
rect 8315 643 8345 695
rect 8397 643 8403 695
rect 5483 630 5736 636
rect 5535 578 5684 630
rect 5483 564 5736 578
rect 5535 512 5684 564
rect 5483 506 5736 512
rect 3018 -63 3287 -21
tri 4571 3 4587 19 se
rect 4587 3 4668 19
tri 4668 3 4702 37 sw
rect 4571 -49 4580 3
rect 4632 -49 4644 3
rect 4696 -49 4702 3
rect 3018 -115 3024 -63
rect 3076 -115 3093 -63
rect 3145 -115 3161 -63
rect 3213 -115 3229 -63
rect 3281 -115 3287 -63
rect 1791 -903 1800 -899
rect 1856 -903 1894 -899
rect 1950 -903 1988 -899
rect 2044 -903 2081 -899
rect 2137 -903 2174 -899
rect 2230 -903 2267 -899
rect 2323 -903 2332 -899
rect 1791 -955 1797 -903
rect 1856 -955 1865 -903
rect 1985 -955 1988 -903
rect 2053 -955 2069 -903
rect 2257 -955 2267 -903
rect 2325 -955 2332 -903
<< via2 >>
rect 7936 1953 7985 1968
rect 7985 1953 7992 1968
rect 8038 1953 8089 1968
rect 8089 1953 8094 1968
rect 7936 1927 7992 1953
rect 8038 1927 8094 1953
rect 7936 1912 7985 1927
rect 7985 1912 7992 1927
rect 8038 1912 8089 1927
rect 8089 1912 8094 1927
rect 8140 1953 8141 1968
rect 8141 1953 8193 1968
rect 8193 1953 8196 1968
rect 8140 1927 8196 1953
rect 8140 1912 8141 1927
rect 8141 1912 8193 1927
rect 8193 1912 8196 1927
rect 8242 1953 8245 1968
rect 8245 1953 8297 1968
rect 8297 1953 8298 1968
rect 8242 1927 8298 1953
rect 8242 1912 8245 1927
rect 8245 1912 8297 1927
rect 8297 1912 8298 1927
rect 8343 1953 8348 1968
rect 8348 1953 8399 1968
rect 8444 1953 8451 1968
rect 8451 1953 8500 1968
rect 8343 1927 8399 1953
rect 8444 1927 8500 1953
rect 8343 1912 8348 1927
rect 8348 1912 8399 1927
rect 8444 1912 8451 1927
rect 8451 1912 8500 1927
rect 7936 793 7985 840
rect 7985 793 7992 840
rect 8035 793 8068 840
rect 8068 793 8091 840
rect 8134 793 8151 840
rect 8151 793 8181 840
rect 8181 793 8190 840
rect 8233 793 8263 840
rect 8263 793 8289 840
rect 8332 793 8345 840
rect 8345 793 8388 840
rect 7936 784 7992 793
rect 8035 784 8091 793
rect 8134 784 8190 793
rect 8233 784 8289 793
rect 8332 784 8388 793
rect 7936 718 7985 760
rect 7985 718 7992 760
rect 8035 718 8068 760
rect 8068 718 8091 760
rect 8134 718 8151 760
rect 8151 718 8181 760
rect 8181 718 8190 760
rect 8233 718 8263 760
rect 8263 718 8289 760
rect 8332 718 8345 760
rect 8345 718 8388 760
rect 7936 704 7992 718
rect 8035 704 8091 718
rect 8134 704 8190 718
rect 8233 704 8289 718
rect 8332 704 8388 718
rect 1800 -903 1856 -899
rect 1894 -903 1950 -899
rect 1988 -903 2044 -899
rect 2081 -903 2137 -899
rect 2174 -903 2230 -899
rect 2267 -903 2323 -899
rect 1800 -955 1849 -903
rect 1849 -955 1856 -903
rect 1894 -955 1917 -903
rect 1917 -955 1933 -903
rect 1933 -955 1950 -903
rect 1988 -955 2001 -903
rect 2001 -955 2044 -903
rect 2081 -955 2121 -903
rect 2121 -955 2137 -903
rect 2174 -955 2189 -903
rect 2189 -955 2205 -903
rect 2205 -955 2230 -903
rect 2267 -955 2273 -903
rect 2273 -955 2323 -903
<< metal3 >>
rect 7931 1968 8505 2010
rect 7931 1912 7936 1968
rect 7992 1912 8038 1968
rect 8094 1912 8140 1968
rect 8196 1912 8242 1968
rect 8298 1912 8343 1968
rect 8399 1912 8444 1968
rect 8500 1912 8505 1968
rect 7931 1870 8505 1912
rect 7931 840 8393 845
rect 7931 784 7936 840
rect 7992 784 8035 840
rect 8091 784 8134 840
rect 8190 784 8233 840
rect 8289 784 8332 840
rect 8388 784 8393 840
rect 7931 760 8393 784
rect 7931 704 7936 760
rect 7992 704 8035 760
rect 8091 704 8134 760
rect 8190 704 8233 760
rect 8289 704 8332 760
rect 8388 704 8393 760
rect 7931 699 8393 704
rect 1795 -899 2328 -894
rect 1795 -955 1800 -899
rect 1856 -955 1894 -899
rect 1950 -955 1988 -899
rect 2044 -955 2081 -899
rect 2137 -955 2174 -899
rect 2230 -955 2267 -899
rect 2323 -955 2328 -899
rect 1795 -960 2328 -955
use sky130_fd_io__com_cclat  sky130_fd_io__com_cclat_0
timestamp 1663361622
transform 1 0 6330 0 1 0
box -133 145 6328 2367
use sky130_fd_io__gpio_dat_ls_1v2  sky130_fd_io__gpio_dat_ls_1v2_0
timestamp 1663361622
transform -1 0 6296 0 -1 2339
box -179 14 3312 2400
use sky130_fd_io__gpio_dat_lsv2  sky130_fd_io__gpio_dat_lsv2_0
timestamp 1663361622
transform 1 0 0 0 -1 2339
box -179 14 3312 2400
use sky130_fd_pr__tpl1__example_55959141808625  sky130_fd_pr__tpl1__example_55959141808625_0
timestamp 1663361622
transform -1 0 6228 0 1 171
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808625  sky130_fd_pr__tpl1__example_55959141808625_1
timestamp 1663361622
transform -1 0 6365 0 1 171
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1663361622
transform -1 0 4689 0 1 -59
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1663361622
transform 1 0 488 0 1 1549
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1663361622
transform -1 0 5903 0 1 1167
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1663361622
transform -1 0 1889 0 1 -49
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1663361622
transform 0 -1 7084 -1 0 1074
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808368  sky130_fd_pr__via_l1m1__example_55959141808368_0
timestamp 1663361622
transform -1 0 12323 0 1 1107
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1663361622
transform 0 -1 6798 -1 0 1030
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1663361622
transform 0 -1 6798 -1 0 1589
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_0
timestamp 1663361622
transform 0 -1 220 -1 0 2004
box 0 0 1 1
<< labels >>
flabel metal2 s 3360 19 3411 49 3 FreeSans 520 0 0 0 OUT
port 1 nsew
flabel metal2 s 2887 19 2933 65 7 FreeSans 300 0 0 0 OE_N
port 2 nsew
flabel metal1 s 7816 1795 7866 1847 3 FreeSans 300 180 0 0 DRVHI_H
port 3 nsew
flabel metal1 s 7493 1715 7545 1767 3 FreeSans 300 180 0 0 DRVLO_H_N
port 4 nsew
flabel metal1 s 12524 2033 12564 2235 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 12433 1875 12473 2005 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 54 1875 94 2005 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s -179 2033 -139 2235 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s -179 884 -139 1086 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 4628 -52 4661 -14 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 7 nsew
flabel metal1 s 5367 93 5434 441 3 FreeSans 520 0 0 0 VPWR_KA
port 8 nsew
flabel locali s 413 1188 448 1234 3 FreeSans 300 0 0 0 OE_H
port 9 nsew
flabel locali s 1048 -30 1110 34 3 FreeSans 520 0 0 0 OD_H
port 10 nsew
flabel comment s 5990 1188 5990 1188 0 FreeSans 300 0 0 0 PU_DIS_H
flabel comment s 6309 1264 6309 1264 0 FreeSans 300 0 0 0 PD_DIS_H
flabel comment s 8460 1325 8460 1325 0 FreeSans 300 0 0 0 PD_DIS_H
flabel comment s 10075 1193 10075 1193 0 FreeSans 300 0 0 0 PD_DIS_H
flabel comment s 6363 1491 6363 1491 0 FreeSans 300 0 0 0 OE_H_N
<< properties >>
string GDS_END 48789786
string GDS_FILE $PDKPATH/libs.ref/gds/sky130_fd_io/sky130_fd_io.gds
string GDS_START 48696232
<< end >>
